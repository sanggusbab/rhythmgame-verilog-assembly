module MemoryControlUnit #(parameter WIDTH = 32,parameter DatamemoryRef = 7788)(counter, PC, Instruction, MemWrite, MemRead, ALUOut, ReadData2,readData,MainGraphic,SingleGraphic,Amplitude,ProgressBar,FrequencyPiezo,LedRGBBright,clockRate);
// if DataAdderss you only need to modify the value of DatamemoryRef
    input[2:0] counter;
    input[WIDTH-1:0] PC;
    input[WIDTH-1:0] ALUOut;
    output reg[WIDTH-1:0] readData;
    output[WIDTH-1:0] Instruction;
    input MemWrite;
    input MemRead;
    input[WIDTH-1:0] ReadData2;

    output[63:0] MainGraphic; // 7368~7375
    output[31:0] SingleGraphic; // 7376~7379
    output[31:0] Amplitude; // 7380~7383
    output[31:0] ProgressBar; // 7384~7387
    output[31:0] FrequencyPiezo; // 7388~7391
    output[31:0] LedRGBBright; // 7392~7395
    output[31:0] clockRate; // 7520~7523
    reg [7:0] Memory [26259:0]; // 8bit per unit Memory - commuticate 32bit
    assign Instruction = {Memory[PC+3],Memory[PC+2],Memory[PC+1],Memory[PC]};

    assign MainGraphic = {Memory[DatamemoryRef+3],Memory[DatamemoryRef+2],Memory[DatamemoryRef+1],Memory[DatamemoryRef],Memory[DatamemoryRef+7],Memory[DatamemoryRef+6],Memory[DatamemoryRef+5],Memory[DatamemoryRef+4]};
    assign SingleGraphic = {Memory[DatamemoryRef+11],Memory[DatamemoryRef+10],Memory[DatamemoryRef+9],Memory[DatamemoryRef+8]};
    assign Amplitude = {Memory[DatamemoryRef+15],Memory[DatamemoryRef+14],Memory[DatamemoryRef+13],Memory[DatamemoryRef+12]};
    assign ProgressBar = {Memory[DatamemoryRef+19],Memory[DatamemoryRef+18],Memory[DatamemoryRef+17],Memory[DatamemoryRef+16]};
    assign FrequencyPiezo = {Memory[DatamemoryRef+23],Memory[DatamemoryRef+22],Memory[DatamemoryRef+21],Memory[DatamemoryRef+20]};
    assign LedRGBBright = {Memory[DatamemoryRef+27],Memory[DatamemoryRef+26],Memory[DatamemoryRef+25],Memory[DatamemoryRef+24]};
    assign clockRate = {Memory[DatamemoryRef+155],Memory[DatamemoryRef+154],Memory[DatamemoryRef+153],Memory[DatamemoryRef+152]};

    always @(counter)begin
        if(counter == 3) begin
            if(MemWrite==1) {Memory[ALUOut+3],Memory[ALUOut+2],Memory[ALUOut+1],Memory[ALUOut]} = ReadData2;
            else if(MemRead) readData = {Memory[ALUOut+3],Memory[ALUOut+2],Memory[ALUOut+1],Memory[ALUOut]};
            else if(~MemRead) readData = ALUOut;
        end
    end
    initial begin
Memory[3] = 8'h00;
Memory[2] = 8'h00;
Memory[1] = 8'h00;
Memory[0] = 8'h93;
Memory[7] = 8'h00;
Memory[6] = 8'h00;
Memory[5] = 8'h01;
Memory[4] = 8'h13;
Memory[11] = 8'h00;
Memory[10] = 8'h00;
Memory[9] = 8'h01;
Memory[8] = 8'h93;
Memory[15] = 8'h00;
Memory[14] = 8'h00;
Memory[13] = 8'h02;
Memory[12] = 8'h13;
Memory[19] = 8'h00;
Memory[18] = 8'h00;
Memory[17] = 8'h02;
Memory[16] = 8'h93;
Memory[23] = 8'h00;
Memory[22] = 8'h00;
Memory[21] = 8'h03;
Memory[20] = 8'h13;
Memory[27] = 8'h00;
Memory[26] = 8'h00;
Memory[25] = 8'h03;
Memory[24] = 8'h93;
Memory[31] = 8'h00;
Memory[30] = 8'h00;
Memory[29] = 8'h04;
Memory[28] = 8'h13;
Memory[35] = 8'h00;
Memory[34] = 8'h00;
Memory[33] = 8'h04;
Memory[32] = 8'h93;
Memory[39] = 8'h00;
Memory[38] = 8'h00;
Memory[37] = 8'h05;
Memory[36] = 8'h13;
Memory[43] = 8'h00;
Memory[42] = 8'h00;
Memory[41] = 8'h05;
Memory[40] = 8'h93;
Memory[47] = 8'h00;
Memory[46] = 8'h00;
Memory[45] = 8'h06;
Memory[44] = 8'h13;
Memory[51] = 8'h00;
Memory[50] = 8'h00;
Memory[49] = 8'h06;
Memory[48] = 8'h93;
Memory[55] = 8'h00;
Memory[54] = 8'h00;
Memory[53] = 8'h07;
Memory[52] = 8'h13;
Memory[59] = 8'h00;
Memory[58] = 8'h00;
Memory[57] = 8'h07;
Memory[56] = 8'h93;
Memory[63] = 8'h00;
Memory[62] = 8'h00;
Memory[61] = 8'h08;
Memory[60] = 8'h13;
Memory[67] = 8'h00;
Memory[66] = 8'h00;
Memory[65] = 8'h08;
Memory[64] = 8'h93;
Memory[71] = 8'h00;
Memory[70] = 8'h00;
Memory[69] = 8'h09;
Memory[68] = 8'h13;
Memory[75] = 8'h00;
Memory[74] = 8'h00;
Memory[73] = 8'h09;
Memory[72] = 8'h93;
Memory[79] = 8'h00;
Memory[78] = 8'h00;
Memory[77] = 8'h0A;
Memory[76] = 8'h13;
Memory[83] = 8'h79;
Memory[82] = 8'hB0;
Memory[81] = 8'h0B;
Memory[80] = 8'h13;
Memory[87] = 8'h00;
Memory[86] = 8'h2B;
Memory[85] = 8'h1B;
Memory[84] = 8'h13;
Memory[91] = 8'h00;
Memory[90] = 8'h00;
Memory[89] = 8'h0B;
Memory[88] = 8'h93;
Memory[95] = 8'h00;
Memory[94] = 8'h10;
Memory[93] = 8'h0C;
Memory[92] = 8'h13;
Memory[99] = 8'h79;
Memory[98] = 8'hF0;
Memory[97] = 8'h0C;
Memory[96] = 8'h93;
Memory[103] = 8'h00;
Memory[102] = 8'h3C;
Memory[101] = 8'h9C;
Memory[100] = 8'h93;
Memory[107] = 8'h21;
Memory[106] = 8'hF0;
Memory[105] = 8'h0D;
Memory[104] = 8'h13;
Memory[111] = 8'h00;
Memory[110] = 8'h5D;
Memory[109] = 8'h1D;
Memory[108] = 8'h13;
Memory[115] = 8'h3E;
Memory[114] = 8'h80;
Memory[113] = 8'h0D;
Memory[112] = 8'h93;
Memory[119] = 8'h00;
Memory[118] = 8'h00;
Memory[117] = 8'h0E;
Memory[116] = 8'h13;
Memory[123] = 8'h00;
Memory[122] = 8'hCC;
Memory[121] = 8'h1B;
Memory[120] = 8'h93;
Memory[127] = 8'h01;
Memory[126] = 8'h3C;
Memory[125] = 8'h1C;
Memory[124] = 8'h13;
Memory[131] = 8'h0A;
Memory[130] = 8'h0B;
Memory[129] = 8'h21;
Memory[128] = 8'h83;
Memory[135] = 8'h0A;
Memory[134] = 8'h4B;
Memory[133] = 8'h22;
Memory[132] = 8'h03;
Memory[139] = 8'h01;
Memory[138] = 8'h10;
Memory[137] = 8'h02;
Memory[136] = 8'h93;
Memory[143] = 8'h00;
Memory[142] = 8'h3B;
Memory[141] = 8'h20;
Memory[140] = 8'h23;
Memory[147] = 8'h00;
Memory[146] = 8'h4B;
Memory[145] = 8'h22;
Memory[144] = 8'h23;
Memory[151] = 8'h00;
Memory[150] = 8'h5B;
Memory[149] = 8'h24;
Memory[148] = 8'h23;
Memory[155] = 8'h00;
Memory[154] = 8'h0B;
Memory[153] = 8'h26;
Memory[152] = 8'h23;
Memory[159] = 8'h01;
Memory[158] = 8'hFF;
Memory[157] = 8'h04;
Memory[156] = 8'h63;
Memory[163] = 8'h11;
Memory[162] = 8'hC0;
Memory[161] = 8'h20;
Memory[160] = 8'h6F;
Memory[167] = 8'h01;
Memory[166] = 8'hDE;
Memory[165] = 8'h14;
Memory[164] = 8'h63;
Memory[171] = 8'hFE;
Memory[170] = 8'h00;
Memory[169] = 8'h0A;
Memory[168] = 8'hE3;
Memory[175] = 8'h00;
Memory[174] = 8'h01;
Memory[173] = 8'h14;
Memory[172] = 8'h63;
Memory[179] = 8'h2C;
Memory[178] = 8'hC0;
Memory[177] = 8'h00;
Memory[176] = 8'h6F;
Memory[183] = 8'h00;
Memory[182] = 8'h10;
Memory[181] = 8'h01;
Memory[180] = 8'h93;
Memory[187] = 8'h00;
Memory[186] = 8'h31;
Memory[185] = 8'h14;
Memory[184] = 8'h63;
Memory[191] = 8'h33;
Memory[190] = 8'h40;
Memory[189] = 8'h00;
Memory[188] = 8'h6F;
Memory[195] = 8'h00;
Memory[194] = 8'h20;
Memory[193] = 8'h01;
Memory[192] = 8'h93;
Memory[199] = 8'h00;
Memory[198] = 8'h31;
Memory[197] = 8'h14;
Memory[196] = 8'h63;
Memory[203] = 8'h38;
Memory[202] = 8'hC0;
Memory[201] = 8'h00;
Memory[200] = 8'h6F;
Memory[207] = 8'h00;
Memory[206] = 8'h30;
Memory[205] = 8'h01;
Memory[204] = 8'h93;
Memory[211] = 8'h00;
Memory[210] = 8'h31;
Memory[209] = 8'h14;
Memory[208] = 8'h63;
Memory[215] = 8'h40;
Memory[214] = 8'h00;
Memory[213] = 8'h00;
Memory[212] = 8'h6F;
Memory[219] = 8'h00;
Memory[218] = 8'h40;
Memory[217] = 8'h01;
Memory[216] = 8'h93;
Memory[223] = 8'h00;
Memory[222] = 8'h31;
Memory[221] = 8'h14;
Memory[220] = 8'h63;
Memory[227] = 8'h48;
Memory[226] = 8'hC0;
Memory[225] = 8'h00;
Memory[224] = 8'h6F;
Memory[231] = 8'h00;
Memory[230] = 8'h50;
Memory[229] = 8'h01;
Memory[228] = 8'h93;
Memory[235] = 8'h00;
Memory[234] = 8'h31;
Memory[233] = 8'h14;
Memory[232] = 8'h63;
Memory[239] = 8'h51;
Memory[238] = 8'h80;
Memory[237] = 8'h00;
Memory[236] = 8'h6F;
Memory[243] = 8'h00;
Memory[242] = 8'h60;
Memory[241] = 8'h01;
Memory[240] = 8'h93;
Memory[247] = 8'h00;
Memory[246] = 8'h31;
Memory[245] = 8'h14;
Memory[244] = 8'h63;
Memory[251] = 8'h5A;
Memory[250] = 8'h40;
Memory[249] = 8'h00;
Memory[248] = 8'h6F;
Memory[255] = 8'h00;
Memory[254] = 8'h70;
Memory[253] = 8'h01;
Memory[252] = 8'h93;
Memory[259] = 8'h00;
Memory[258] = 8'h31;
Memory[257] = 8'h14;
Memory[256] = 8'h63;
Memory[263] = 8'h63;
Memory[262] = 8'h00;
Memory[261] = 8'h00;
Memory[260] = 8'h6F;
Memory[267] = 8'h00;
Memory[266] = 8'h80;
Memory[265] = 8'h01;
Memory[264] = 8'h93;
Memory[271] = 8'h00;
Memory[270] = 8'h31;
Memory[269] = 8'h14;
Memory[268] = 8'h63;
Memory[275] = 8'h6A;
Memory[274] = 8'h80;
Memory[273] = 8'h00;
Memory[272] = 8'h6F;
Memory[279] = 8'h00;
Memory[278] = 8'h90;
Memory[277] = 8'h01;
Memory[276] = 8'h93;
Memory[283] = 8'h00;
Memory[282] = 8'h31;
Memory[281] = 8'h14;
Memory[280] = 8'h63;
Memory[287] = 8'h71;
Memory[286] = 8'h80;
Memory[285] = 8'h00;
Memory[284] = 8'h6F;
Memory[291] = 8'h00;
Memory[290] = 8'hA0;
Memory[289] = 8'h01;
Memory[288] = 8'h93;
Memory[295] = 8'h00;
Memory[294] = 8'h31;
Memory[293] = 8'h14;
Memory[292] = 8'h63;
Memory[299] = 8'h79;
Memory[298] = 8'hC0;
Memory[297] = 8'h00;
Memory[296] = 8'h6F;
Memory[303] = 8'h00;
Memory[302] = 8'hB0;
Memory[301] = 8'h01;
Memory[300] = 8'h93;
Memory[307] = 8'h00;
Memory[306] = 8'h31;
Memory[305] = 8'h14;
Memory[304] = 8'h63;
Memory[311] = 8'h08;
Memory[310] = 8'h90;
Memory[309] = 8'h00;
Memory[308] = 8'h6F;
Memory[315] = 8'h00;
Memory[314] = 8'hC0;
Memory[313] = 8'h01;
Memory[312] = 8'h93;
Memory[319] = 8'h00;
Memory[318] = 8'h31;
Memory[317] = 8'h14;
Memory[316] = 8'h63;
Memory[323] = 8'h18;
Memory[322] = 8'h90;
Memory[321] = 8'h00;
Memory[320] = 8'h6F;
Memory[327] = 8'h00;
Memory[326] = 8'hD0;
Memory[325] = 8'h01;
Memory[324] = 8'h93;
Memory[331] = 8'h00;
Memory[330] = 8'h31;
Memory[329] = 8'h14;
Memory[328] = 8'h63;
Memory[335] = 8'h28;
Memory[334] = 8'h90;
Memory[333] = 8'h00;
Memory[332] = 8'h6F;
Memory[339] = 8'h01;
Memory[338] = 8'h30;
Memory[337] = 8'h01;
Memory[336] = 8'h93;
Memory[343] = 8'h00;
Memory[342] = 8'h31;
Memory[341] = 8'h14;
Memory[340] = 8'h63;
Memory[347] = 8'h37;
Memory[346] = 8'h50;
Memory[345] = 8'h00;
Memory[344] = 8'h6F;
Memory[351] = 8'h01;
Memory[350] = 8'h40;
Memory[349] = 8'h01;
Memory[348] = 8'h93;
Memory[355] = 8'h00;
Memory[354] = 8'h31;
Memory[353] = 8'h14;
Memory[352] = 8'h63;
Memory[359] = 8'h3F;
Memory[358] = 8'hD0;
Memory[357] = 8'h00;
Memory[356] = 8'h6F;
Memory[363] = 8'h01;
Memory[362] = 8'h50;
Memory[361] = 8'h01;
Memory[360] = 8'h93;
Memory[367] = 8'h00;
Memory[366] = 8'h31;
Memory[365] = 8'h14;
Memory[364] = 8'h63;
Memory[371] = 8'h46;
Memory[370] = 8'h90;
Memory[369] = 8'h00;
Memory[368] = 8'h6F;
Memory[375] = 8'h01;
Memory[374] = 8'h60;
Memory[373] = 8'h01;
Memory[372] = 8'h93;
Memory[379] = 8'h00;
Memory[378] = 8'h31;
Memory[377] = 8'h14;
Memory[376] = 8'h63;
Memory[383] = 8'h4E;
Memory[382] = 8'h90;
Memory[381] = 8'h00;
Memory[380] = 8'h6F;
Memory[387] = 8'h01;
Memory[386] = 8'h70;
Memory[385] = 8'h01;
Memory[384] = 8'h93;
Memory[391] = 8'h00;
Memory[390] = 8'h31;
Memory[389] = 8'h14;
Memory[388] = 8'h63;
Memory[395] = 8'h56;
Memory[394] = 8'h90;
Memory[393] = 8'h00;
Memory[392] = 8'h6F;
Memory[399] = 8'h01;
Memory[398] = 8'h80;
Memory[397] = 8'h01;
Memory[396] = 8'h93;
Memory[403] = 8'h00;
Memory[402] = 8'h31;
Memory[401] = 8'h14;
Memory[400] = 8'h63;
Memory[407] = 8'h5E;
Memory[406] = 8'h90;
Memory[405] = 8'h00;
Memory[404] = 8'h6F;
Memory[411] = 8'h01;
Memory[410] = 8'h90;
Memory[409] = 8'h01;
Memory[408] = 8'h93;
Memory[415] = 8'h00;
Memory[414] = 8'h31;
Memory[413] = 8'h14;
Memory[412] = 8'h63;
Memory[419] = 8'h66;
Memory[418] = 8'h90;
Memory[417] = 8'h00;
Memory[416] = 8'h6F;
Memory[423] = 8'h01;
Memory[422] = 8'hA0;
Memory[421] = 8'h01;
Memory[420] = 8'h93;
Memory[427] = 8'h00;
Memory[426] = 8'h31;
Memory[425] = 8'h14;
Memory[424] = 8'h63;
Memory[431] = 8'h6E;
Memory[430] = 8'h90;
Memory[429] = 8'h00;
Memory[428] = 8'h6F;
Memory[435] = 8'h01;
Memory[434] = 8'hB0;
Memory[433] = 8'h01;
Memory[432] = 8'h93;
Memory[439] = 8'h00;
Memory[438] = 8'h31;
Memory[437] = 8'h14;
Memory[436] = 8'h63;
Memory[443] = 8'h76;
Memory[442] = 8'h90;
Memory[441] = 8'h00;
Memory[440] = 8'h6F;
Memory[447] = 8'h01;
Memory[446] = 8'hC0;
Memory[445] = 8'h01;
Memory[444] = 8'h93;
Memory[451] = 8'h00;
Memory[450] = 8'h31;
Memory[449] = 8'h14;
Memory[448] = 8'h63;
Memory[455] = 8'h7D;
Memory[454] = 8'h50;
Memory[453] = 8'h00;
Memory[452] = 8'h6F;
Memory[459] = 8'h01;
Memory[458] = 8'hD0;
Memory[457] = 8'h01;
Memory[456] = 8'h93;
Memory[463] = 8'h00;
Memory[462] = 8'h31;
Memory[461] = 8'h14;
Memory[460] = 8'h63;
Memory[467] = 8'h04;
Memory[466] = 8'h80;
Memory[465] = 8'h10;
Memory[464] = 8'h6F;
Memory[471] = 8'h01;
Memory[470] = 8'hE0;
Memory[469] = 8'h01;
Memory[468] = 8'h93;
Memory[475] = 8'h00;
Memory[474] = 8'h31;
Memory[473] = 8'h14;
Memory[472] = 8'h63;
Memory[479] = 8'h0D;
Memory[478] = 8'h00;
Memory[477] = 8'h10;
Memory[476] = 8'h6F;
Memory[483] = 8'h01;
Memory[482] = 8'hF0;
Memory[481] = 8'h01;
Memory[480] = 8'h93;
Memory[487] = 8'h00;
Memory[486] = 8'h31;
Memory[485] = 8'h14;
Memory[484] = 8'h63;
Memory[491] = 8'h32;
Memory[490] = 8'h40;
Memory[489] = 8'h10;
Memory[488] = 8'h6F;
Memory[495] = 8'h02;
Memory[494] = 8'h00;
Memory[493] = 8'h01;
Memory[492] = 8'h93;
Memory[499] = 8'h00;
Memory[498] = 8'h31;
Memory[497] = 8'h14;
Memory[496] = 8'h63;
Memory[503] = 8'h3A;
Memory[502] = 8'hC0;
Memory[501] = 8'h10;
Memory[500] = 8'h6F;
Memory[507] = 8'h02;
Memory[506] = 8'h10;
Memory[505] = 8'h01;
Memory[504] = 8'h93;
Memory[511] = 8'h00;
Memory[510] = 8'h31;
Memory[509] = 8'h14;
Memory[508] = 8'h63;
Memory[515] = 8'h60;
Memory[514] = 8'h00;
Memory[513] = 8'h10;
Memory[512] = 8'h6F;
Memory[519] = 8'h02;
Memory[518] = 8'h50;
Memory[517] = 8'h01;
Memory[516] = 8'h93;
Memory[523] = 8'h00;
Memory[522] = 8'h31;
Memory[521] = 8'h14;
Memory[520] = 8'h63;
Memory[527] = 8'h67;
Memory[526] = 8'h40;
Memory[525] = 8'h10;
Memory[524] = 8'h6F;
Memory[531] = 8'h02;
Memory[530] = 8'h60;
Memory[529] = 8'h01;
Memory[528] = 8'h93;
Memory[535] = 8'h00;
Memory[534] = 8'h31;
Memory[533] = 8'h14;
Memory[532] = 8'h63;
Memory[539] = 8'h6F;
Memory[538] = 8'hC0;
Memory[537] = 8'h10;
Memory[536] = 8'h6F;
Memory[543] = 8'h02;
Memory[542] = 8'h70;
Memory[541] = 8'h01;
Memory[540] = 8'h93;
Memory[547] = 8'h00;
Memory[546] = 8'h31;
Memory[545] = 8'h14;
Memory[544] = 8'h63;
Memory[551] = 8'h78;
Memory[550] = 8'h40;
Memory[549] = 8'h10;
Memory[548] = 8'h6F;
Memory[555] = 8'h02;
Memory[554] = 8'h80;
Memory[553] = 8'h01;
Memory[552] = 8'h93;
Memory[559] = 8'h00;
Memory[558] = 8'h31;
Memory[557] = 8'h14;
Memory[556] = 8'h63;
Memory[563] = 8'h01;
Memory[562] = 8'hD0;
Memory[561] = 8'h10;
Memory[560] = 8'h6F;
Memory[567] = 8'h02;
Memory[566] = 8'h90;
Memory[565] = 8'h01;
Memory[564] = 8'h93;
Memory[571] = 8'h00;
Memory[570] = 8'h31;
Memory[569] = 8'h14;
Memory[568] = 8'h63;
Memory[575] = 8'h0B;
Memory[574] = 8'h50;
Memory[573] = 8'h10;
Memory[572] = 8'h6F;
Memory[579] = 8'h02;
Memory[578] = 8'hA0;
Memory[577] = 8'h01;
Memory[576] = 8'h93;
Memory[583] = 8'h00;
Memory[582] = 8'h31;
Memory[581] = 8'h14;
Memory[580] = 8'h63;
Memory[587] = 8'h14;
Memory[586] = 8'hD0;
Memory[585] = 8'h10;
Memory[584] = 8'h6F;
Memory[591] = 8'h02;
Memory[590] = 8'hB0;
Memory[589] = 8'h01;
Memory[588] = 8'h93;
Memory[595] = 8'h00;
Memory[594] = 8'h31;
Memory[593] = 8'h14;
Memory[592] = 8'h63;
Memory[599] = 8'h1E;
Memory[598] = 8'h50;
Memory[597] = 8'h10;
Memory[596] = 8'h6F;
Memory[603] = 8'h02;
Memory[602] = 8'hE0;
Memory[601] = 8'h01;
Memory[600] = 8'h93;
Memory[607] = 8'h00;
Memory[606] = 8'h31;
Memory[605] = 8'h14;
Memory[604] = 8'h63;
Memory[611] = 8'h23;
Memory[610] = 8'h10;
Memory[609] = 8'h10;
Memory[608] = 8'h6F;
Memory[615] = 8'h02;
Memory[614] = 8'hF0;
Memory[613] = 8'h01;
Memory[612] = 8'h93;
Memory[619] = 8'h00;
Memory[618] = 8'h31;
Memory[617] = 8'h14;
Memory[616] = 8'h63;
Memory[623] = 8'h2C;
Memory[622] = 8'h90;
Memory[621] = 8'h10;
Memory[620] = 8'h6F;
Memory[627] = 8'h03;
Memory[626] = 8'h00;
Memory[625] = 8'h01;
Memory[624] = 8'h93;
Memory[631] = 8'h00;
Memory[630] = 8'h31;
Memory[629] = 8'h14;
Memory[628] = 8'h63;
Memory[635] = 8'h35;
Memory[634] = 8'hD0;
Memory[633] = 8'h10;
Memory[632] = 8'h6F;
Memory[639] = 8'h03;
Memory[638] = 8'h10;
Memory[637] = 8'h01;
Memory[636] = 8'h93;
Memory[643] = 8'h00;
Memory[642] = 8'h31;
Memory[641] = 8'h14;
Memory[640] = 8'h63;
Memory[647] = 8'h40;
Memory[646] = 8'hD0;
Memory[645] = 8'h10;
Memory[644] = 8'h6F;
Memory[651] = 8'h03;
Memory[650] = 8'h20;
Memory[649] = 8'h01;
Memory[648] = 8'h93;
Memory[655] = 8'h00;
Memory[654] = 8'h31;
Memory[653] = 8'h14;
Memory[652] = 8'h63;
Memory[659] = 8'h4A;
Memory[658] = 8'h10;
Memory[657] = 8'h10;
Memory[656] = 8'h6F;
Memory[663] = 8'h03;
Memory[662] = 8'h40;
Memory[661] = 8'h01;
Memory[660] = 8'h93;
Memory[667] = 8'h00;
Memory[666] = 8'h31;
Memory[665] = 8'h14;
Memory[664] = 8'h63;
Memory[671] = 8'h50;
Memory[670] = 8'h90;
Memory[669] = 8'h10;
Memory[668] = 8'h6F;
Memory[675] = 8'h03;
Memory[674] = 8'h60;
Memory[673] = 8'h01;
Memory[672] = 8'h93;
Memory[679] = 8'h00;
Memory[678] = 8'h31;
Memory[677] = 8'h14;
Memory[676] = 8'h63;
Memory[683] = 8'h55;
Memory[682] = 8'hD0;
Memory[681] = 8'h10;
Memory[680] = 8'h6F;
Memory[687] = 8'h03;
Memory[686] = 8'h70;
Memory[685] = 8'h01;
Memory[684] = 8'h93;
Memory[691] = 8'h00;
Memory[690] = 8'h31;
Memory[689] = 8'h14;
Memory[688] = 8'h63;
Memory[695] = 8'h5B;
Memory[694] = 8'h10;
Memory[693] = 8'h10;
Memory[692] = 8'h6F;
Memory[699] = 8'h03;
Memory[698] = 8'h80;
Memory[697] = 8'h01;
Memory[696] = 8'h93;
Memory[703] = 8'h00;
Memory[702] = 8'h31;
Memory[701] = 8'h14;
Memory[700] = 8'h63;
Memory[707] = 8'h0D;
Memory[706] = 8'h00;
Memory[705] = 8'h20;
Memory[704] = 8'h6F;
Memory[711] = 8'h00;
Memory[710] = 8'h0E;
Memory[709] = 8'h8E;
Memory[708] = 8'h13;
Memory[715] = 8'hDC;
Memory[714] = 8'h00;
Memory[713] = 8'h0A;
Memory[712] = 8'hE3;
Memory[719] = 8'h00;
Memory[718] = 8'h00;
Memory[717] = 8'h01;
Memory[716] = 8'h13;
Memory[723] = 8'h0A;
Memory[722] = 8'h0B;
Memory[721] = 8'h21;
Memory[720] = 8'h83;
Memory[727] = 8'h0A;
Memory[726] = 8'h4B;
Memory[725] = 8'h22;
Memory[724] = 8'h03;
Memory[731] = 8'h01;
Memory[730] = 8'h10;
Memory[729] = 8'h02;
Memory[728] = 8'h93;
Memory[735] = 8'h00;
Memory[734] = 8'h3B;
Memory[733] = 8'h20;
Memory[732] = 8'h23;
Memory[739] = 8'h00;
Memory[738] = 8'h4B;
Memory[737] = 8'h22;
Memory[736] = 8'h23;
Memory[743] = 8'h00;
Memory[742] = 8'h5B;
Memory[741] = 8'h24;
Memory[740] = 8'h23;
Memory[747] = 8'h00;
Memory[746] = 8'h0B;
Memory[745] = 8'h26;
Memory[744] = 8'h23;
Memory[751] = 8'h01;
Memory[750] = 8'hDE;
Memory[749] = 8'h14;
Memory[748] = 8'h63;
Memory[755] = 8'h09;
Memory[754] = 8'hC0;
Memory[753] = 8'h00;
Memory[752] = 8'h6F;
Memory[759] = 8'h01;
Memory[758] = 8'hDE;
Memory[757] = 8'h42;
Memory[756] = 8'h33;
Memory[763] = 8'h01;
Memory[762] = 8'h82;
Memory[761] = 8'h71;
Memory[760] = 8'hB3;
Memory[767] = 8'h01;
Memory[766] = 8'hD1;
Memory[765] = 8'hF1;
Memory[764] = 8'hB3;
Memory[771] = 8'h00;
Memory[770] = 8'h01;
Memory[769] = 8'h84;
Memory[768] = 8'h63;
Memory[775] = 8'h0D;
Memory[774] = 8'h00;
Memory[773] = 8'h20;
Memory[772] = 8'h6F;
Memory[779] = 8'hFF;
Memory[778] = 8'hF2;
Memory[777] = 8'h71;
Memory[776] = 8'h93;
Memory[783] = 8'h01;
Memory[782] = 8'hD1;
Memory[781] = 8'hF1;
Memory[780] = 8'hB3;
Memory[787] = 8'hFA;
Memory[786] = 8'h01;
Memory[785] = 8'h8A;
Memory[784] = 8'hE3;
Memory[791] = 8'h0A;
Memory[790] = 8'h8B;
Memory[789] = 8'h21;
Memory[788] = 8'h83;
Memory[795] = 8'h0A;
Memory[794] = 8'hCB;
Memory[793] = 8'h22;
Memory[792] = 8'h03;
Memory[799] = 8'h29;
Memory[798] = 8'h8B;
Memory[797] = 8'h22;
Memory[796] = 8'h83;
Memory[803] = 8'h00;
Memory[802] = 8'h3B;
Memory[801] = 8'h20;
Memory[800] = 8'h23;
Memory[807] = 8'h00;
Memory[806] = 8'h4B;
Memory[805] = 8'h22;
Memory[804] = 8'h23;
Memory[811] = 8'h00;
Memory[810] = 8'h5B;
Memory[809] = 8'h24;
Memory[808] = 8'h23;
Memory[815] = 8'h00;
Memory[814] = 8'h10;
Memory[813] = 8'h01;
Memory[812] = 8'h13;
Memory[819] = 8'h2C;
Memory[818] = 8'h40;
Memory[817] = 8'h00;
Memory[816] = 8'h6F;
Memory[823] = 8'h00;
Memory[822] = 8'h10;
Memory[821] = 8'h01;
Memory[820] = 8'h13;
Memory[827] = 8'h0A;
Memory[826] = 8'h8B;
Memory[825] = 8'h21;
Memory[824] = 8'h83;
Memory[831] = 8'h0A;
Memory[830] = 8'hCB;
Memory[829] = 8'h22;
Memory[828] = 8'h03;
Memory[835] = 8'h29;
Memory[834] = 8'h8B;
Memory[833] = 8'h22;
Memory[832] = 8'h83;
Memory[839] = 8'h00;
Memory[838] = 8'h3B;
Memory[837] = 8'h20;
Memory[836] = 8'h23;
Memory[843] = 8'h00;
Memory[842] = 8'h4B;
Memory[841] = 8'h22;
Memory[840] = 8'h23;
Memory[847] = 8'h00;
Memory[846] = 8'h5B;
Memory[845] = 8'h24;
Memory[844] = 8'h23;
Memory[851] = 8'h01;
Memory[850] = 8'hDE;
Memory[849] = 8'h14;
Memory[848] = 8'h63;
Memory[855] = 8'h09;
Memory[854] = 8'hC0;
Memory[853] = 8'h00;
Memory[852] = 8'h6F;
Memory[859] = 8'h01;
Memory[858] = 8'hDE;
Memory[857] = 8'h42;
Memory[856] = 8'h33;
Memory[863] = 8'h01;
Memory[862] = 8'h82;
Memory[861] = 8'h71;
Memory[860] = 8'hB3;
Memory[867] = 8'h01;
Memory[866] = 8'hD1;
Memory[865] = 8'hF1;
Memory[864] = 8'hB3;
Memory[871] = 8'h00;
Memory[870] = 8'h01;
Memory[869] = 8'h84;
Memory[868] = 8'h63;
Memory[875] = 8'h0D;
Memory[874] = 8'h00;
Memory[873] = 8'h20;
Memory[872] = 8'h6F;
Memory[879] = 8'hFF;
Memory[878] = 8'hF2;
Memory[877] = 8'h71;
Memory[876] = 8'h93;
Memory[883] = 8'h01;
Memory[882] = 8'hD1;
Memory[881] = 8'hF1;
Memory[880] = 8'hB3;
Memory[887] = 8'hF4;
Memory[886] = 8'h01;
Memory[885] = 8'h88;
Memory[884] = 8'hE3;
Memory[891] = 8'h0B;
Memory[890] = 8'h0B;
Memory[889] = 8'h21;
Memory[888] = 8'h83;
Memory[895] = 8'h0B;
Memory[894] = 8'h4B;
Memory[893] = 8'h22;
Memory[892] = 8'h03;
Memory[899] = 8'h00;
Memory[898] = 8'h3B;
Memory[897] = 8'h20;
Memory[896] = 8'h23;
Memory[903] = 8'h00;
Memory[902] = 8'h4B;
Memory[901] = 8'h22;
Memory[900] = 8'h23;
Memory[907] = 8'h38;
Memory[906] = 8'hC0;
Memory[905] = 8'h00;
Memory[904] = 8'h6F;
Memory[911] = 8'h00;
Memory[910] = 8'h20;
Memory[909] = 8'h01;
Memory[908] = 8'h13;
Memory[915] = 8'h0B;
Memory[914] = 8'h0B;
Memory[913] = 8'h21;
Memory[912] = 8'h83;
Memory[919] = 8'h0B;
Memory[918] = 8'h4B;
Memory[917] = 8'h22;
Memory[916] = 8'h03;
Memory[923] = 8'h00;
Memory[922] = 8'h3B;
Memory[921] = 8'h20;
Memory[920] = 8'h23;
Memory[927] = 8'h00;
Memory[926] = 8'h4B;
Memory[925] = 8'h22;
Memory[924] = 8'h23;
Memory[931] = 8'h01;
Memory[930] = 8'hDE;
Memory[929] = 8'h14;
Memory[928] = 8'h63;
Memory[935] = 8'h09;
Memory[934] = 8'hC0;
Memory[933] = 8'h00;
Memory[932] = 8'h6F;
Memory[939] = 8'h01;
Memory[938] = 8'hDE;
Memory[937] = 8'h42;
Memory[936] = 8'h33;
Memory[943] = 8'h01;
Memory[942] = 8'h82;
Memory[941] = 8'h71;
Memory[940] = 8'hB3;
Memory[947] = 8'h01;
Memory[946] = 8'hD1;
Memory[945] = 8'hF1;
Memory[944] = 8'hB3;
Memory[951] = 8'h00;
Memory[950] = 8'h01;
Memory[949] = 8'h84;
Memory[948] = 8'h63;
Memory[955] = 8'h0D;
Memory[954] = 8'h00;
Memory[953] = 8'h20;
Memory[952] = 8'h6F;
Memory[959] = 8'hFF;
Memory[958] = 8'hF2;
Memory[957] = 8'h71;
Memory[956] = 8'h93;
Memory[963] = 8'h01;
Memory[962] = 8'hD1;
Memory[961] = 8'hF1;
Memory[960] = 8'hB3;
Memory[967] = 8'hF0;
Memory[966] = 8'h01;
Memory[965] = 8'h80;
Memory[964] = 8'hE3;
Memory[971] = 8'h01;
Memory[970] = 8'h01;
Memory[969] = 8'hF2;
Memory[968] = 8'h13;
Memory[975] = 8'h00;
Memory[974] = 8'h02;
Memory[973] = 8'h18;
Memory[972] = 8'h63;
Memory[979] = 8'h00;
Memory[978] = 8'h41;
Memory[977] = 8'hF2;
Memory[976] = 8'h13;
Memory[983] = 8'h00;
Memory[982] = 8'h02;
Memory[981] = 8'h1A;
Memory[980] = 8'h63;
Memory[987] = 8'h2C;
Memory[986] = 8'h40;
Memory[985] = 8'h00;
Memory[984] = 8'h6F;
Memory[991] = 8'h00;
Memory[990] = 8'h30;
Memory[989] = 8'h01;
Memory[988] = 8'h13;
Memory[995] = 8'h00;
Memory[994] = 8'h0E;
Memory[993] = 8'h8E;
Memory[992] = 8'h13;
Memory[999] = 8'h00;
Memory[998] = 8'h00;
Memory[997] = 8'h0E;
Memory[996] = 8'h63;
Memory[1003] = 8'h01;
Memory[1002] = 8'hB0;
Memory[1001] = 8'h01;
Memory[1000] = 8'hB3;
Memory[1007] = 8'h03;
Memory[1006] = 8'hB1;
Memory[1005] = 8'h81;
Memory[1004] = 8'hB3;
Memory[1011] = 8'h08;
Memory[1010] = 8'h3B;
Memory[1009] = 8'h2C;
Memory[1008] = 8'h23;
Memory[1015] = 8'h00;
Memory[1014] = 8'h80;
Memory[1013] = 8'h01;
Memory[1012] = 8'h13;
Memory[1019] = 8'h00;
Memory[1018] = 8'h0E;
Memory[1017] = 8'h8E;
Memory[1016] = 8'h13;
Memory[1023] = 8'h2A;
Memory[1022] = 8'h00;
Memory[1021] = 8'h06;
Memory[1020] = 8'h63;
Memory[1027] = 8'h00;
Memory[1026] = 8'h30;
Memory[1025] = 8'h01;
Memory[1024] = 8'h13;
Memory[1031] = 8'h0B;
Memory[1030] = 8'h8B;
Memory[1029] = 8'h21;
Memory[1028] = 8'h83;
Memory[1035] = 8'h0B;
Memory[1034] = 8'hCB;
Memory[1033] = 8'h22;
Memory[1032] = 8'h03;
Memory[1039] = 8'h00;
Memory[1038] = 8'h3B;
Memory[1037] = 8'h20;
Memory[1036] = 8'h23;
Memory[1043] = 8'h00;
Memory[1042] = 8'h4B;
Memory[1041] = 8'h22;
Memory[1040] = 8'h23;
Memory[1047] = 8'h01;
Memory[1046] = 8'hDE;
Memory[1045] = 8'h14;
Memory[1044] = 8'h63;
Memory[1051] = 8'h09;
Memory[1050] = 8'hC0;
Memory[1049] = 8'h00;
Memory[1048] = 8'h6F;
Memory[1055] = 8'h01;
Memory[1054] = 8'hDE;
Memory[1053] = 8'h42;
Memory[1052] = 8'h33;
Memory[1059] = 8'h01;
Memory[1058] = 8'h82;
Memory[1057] = 8'h71;
Memory[1056] = 8'hB3;
Memory[1063] = 8'h01;
Memory[1062] = 8'hD1;
Memory[1061] = 8'hF1;
Memory[1060] = 8'hB3;
Memory[1067] = 8'h00;
Memory[1066] = 8'h01;
Memory[1065] = 8'h84;
Memory[1064] = 8'h63;
Memory[1071] = 8'h0D;
Memory[1070] = 8'h00;
Memory[1069] = 8'h20;
Memory[1068] = 8'h6F;
Memory[1075] = 8'hFF;
Memory[1074] = 8'hF2;
Memory[1073] = 8'h71;
Memory[1072] = 8'h93;
Memory[1079] = 8'h01;
Memory[1078] = 8'hD1;
Memory[1077] = 8'hF1;
Memory[1076] = 8'hB3;
Memory[1083] = 8'hE8;
Memory[1082] = 8'h01;
Memory[1081] = 8'h86;
Memory[1080] = 8'hE3;
Memory[1087] = 8'h40;
Memory[1086] = 8'h01;
Memory[1085] = 8'hF2;
Memory[1084] = 8'h13;
Memory[1091] = 8'h00;
Memory[1090] = 8'h02;
Memory[1089] = 8'h1C;
Memory[1088] = 8'h63;
Memory[1095] = 8'h01;
Memory[1094] = 8'h01;
Memory[1093] = 8'hF2;
Memory[1092] = 8'h13;
Memory[1099] = 8'h00;
Memory[1098] = 8'h02;
Memory[1097] = 8'h1E;
Memory[1096] = 8'h63;
Memory[1103] = 8'h00;
Memory[1102] = 8'h41;
Memory[1101] = 8'hF2;
Memory[1100] = 8'h13;
Memory[1107] = 8'h02;
Memory[1106] = 8'h02;
Memory[1105] = 8'h10;
Memory[1104] = 8'h63;
Memory[1111] = 8'h2C;
Memory[1110] = 8'h40;
Memory[1109] = 8'h00;
Memory[1108] = 8'h6F;
Memory[1115] = 8'h00;
Memory[1114] = 8'h20;
Memory[1113] = 8'h01;
Memory[1112] = 8'h13;
Memory[1119] = 8'h00;
Memory[1118] = 8'h0E;
Memory[1117] = 8'h8E;
Memory[1116] = 8'h13;
Memory[1123] = 8'hF2;
Memory[1122] = 8'h00;
Memory[1121] = 8'h06;
Memory[1120] = 8'hE3;
Memory[1127] = 8'h00;
Memory[1126] = 8'h40;
Memory[1125] = 8'h01;
Memory[1124] = 8'h13;
Memory[1131] = 8'h00;
Memory[1130] = 8'h0E;
Memory[1129] = 8'h8E;
Memory[1128] = 8'h13;
Memory[1135] = 8'h02;
Memory[1134] = 8'h00;
Memory[1133] = 8'h00;
Memory[1132] = 8'h63;
Memory[1139] = 8'h00;
Memory[1138] = 8'hA0;
Memory[1137] = 8'h01;
Memory[1136] = 8'h93;
Memory[1143] = 8'h03;
Memory[1142] = 8'hB1;
Memory[1141] = 8'h81;
Memory[1140] = 8'hB3;
Memory[1147] = 8'h03;
Memory[1146] = 8'hB1;
Memory[1145] = 8'h81;
Memory[1144] = 8'hB3;
Memory[1151] = 8'h08;
Memory[1150] = 8'h3B;
Memory[1149] = 8'h2C;
Memory[1148] = 8'h23;
Memory[1155] = 8'h00;
Memory[1154] = 8'h80;
Memory[1153] = 8'h01;
Memory[1152] = 8'h13;
Memory[1159] = 8'h00;
Memory[1158] = 8'h0E;
Memory[1157] = 8'h8E;
Memory[1156] = 8'h13;
Memory[1163] = 8'h22;
Memory[1162] = 8'h00;
Memory[1161] = 8'h00;
Memory[1160] = 8'h63;
Memory[1167] = 8'h00;
Memory[1166] = 8'h40;
Memory[1165] = 8'h01;
Memory[1164] = 8'h13;
Memory[1171] = 8'h0C;
Memory[1170] = 8'h0B;
Memory[1169] = 8'h21;
Memory[1168] = 8'h83;
Memory[1175] = 8'h0C;
Memory[1174] = 8'h4B;
Memory[1173] = 8'h22;
Memory[1172] = 8'h03;
Memory[1179] = 8'h00;
Memory[1178] = 8'h3B;
Memory[1177] = 8'h20;
Memory[1176] = 8'h23;
Memory[1183] = 8'h00;
Memory[1182] = 8'h4B;
Memory[1181] = 8'h22;
Memory[1180] = 8'h23;
Memory[1187] = 8'h01;
Memory[1186] = 8'hDE;
Memory[1185] = 8'h14;
Memory[1184] = 8'h63;
Memory[1191] = 8'h09;
Memory[1190] = 8'hC0;
Memory[1189] = 8'h00;
Memory[1188] = 8'h6F;
Memory[1195] = 8'h01;
Memory[1194] = 8'hDE;
Memory[1193] = 8'h42;
Memory[1192] = 8'h33;
Memory[1199] = 8'h01;
Memory[1198] = 8'h82;
Memory[1197] = 8'h71;
Memory[1196] = 8'hB3;
Memory[1203] = 8'h01;
Memory[1202] = 8'hD1;
Memory[1201] = 8'hF1;
Memory[1200] = 8'hB3;
Memory[1207] = 8'h00;
Memory[1206] = 8'h01;
Memory[1205] = 8'h84;
Memory[1204] = 8'h63;
Memory[1211] = 8'h0D;
Memory[1210] = 8'h00;
Memory[1209] = 8'h20;
Memory[1208] = 8'h6F;
Memory[1215] = 8'hFF;
Memory[1214] = 8'hF2;
Memory[1213] = 8'h71;
Memory[1212] = 8'h93;
Memory[1219] = 8'h01;
Memory[1218] = 8'hD1;
Memory[1217] = 8'hF1;
Memory[1216] = 8'hB3;
Memory[1223] = 8'hE0;
Memory[1222] = 8'h01;
Memory[1221] = 8'h80;
Memory[1220] = 8'hE3;
Memory[1227] = 8'h40;
Memory[1226] = 8'h01;
Memory[1225] = 8'hF2;
Memory[1224] = 8'h13;
Memory[1231] = 8'h00;
Memory[1230] = 8'h02;
Memory[1229] = 8'h1C;
Memory[1228] = 8'h63;
Memory[1235] = 8'h01;
Memory[1234] = 8'h01;
Memory[1233] = 8'hF2;
Memory[1232] = 8'h13;
Memory[1239] = 8'h00;
Memory[1238] = 8'h02;
Memory[1237] = 8'h1E;
Memory[1236] = 8'h63;
Memory[1243] = 8'h00;
Memory[1242] = 8'h41;
Memory[1241] = 8'hF2;
Memory[1240] = 8'h13;
Memory[1247] = 8'h02;
Memory[1246] = 8'h02;
Memory[1245] = 8'h10;
Memory[1244] = 8'h63;
Memory[1251] = 8'h2C;
Memory[1250] = 8'h40;
Memory[1249] = 8'h00;
Memory[1248] = 8'h6F;
Memory[1255] = 8'h00;
Memory[1254] = 8'h30;
Memory[1253] = 8'h01;
Memory[1252] = 8'h13;
Memory[1259] = 8'h00;
Memory[1258] = 8'h0E;
Memory[1257] = 8'h8E;
Memory[1256] = 8'h13;
Memory[1263] = 8'hF0;
Memory[1262] = 8'h00;
Memory[1261] = 8'h0A;
Memory[1260] = 8'hE3;
Memory[1267] = 8'h00;
Memory[1266] = 8'h50;
Memory[1265] = 8'h01;
Memory[1264] = 8'h13;
Memory[1271] = 8'h00;
Memory[1270] = 8'h0E;
Memory[1269] = 8'h8E;
Memory[1268] = 8'h13;
Memory[1275] = 8'h02;
Memory[1274] = 8'h00;
Memory[1273] = 8'h00;
Memory[1272] = 8'h63;
Memory[1279] = 8'h03;
Memory[1278] = 8'h20;
Memory[1277] = 8'h01;
Memory[1276] = 8'h93;
Memory[1283] = 8'h03;
Memory[1282] = 8'hB1;
Memory[1281] = 8'h81;
Memory[1280] = 8'hB3;
Memory[1287] = 8'h03;
Memory[1286] = 8'hB1;
Memory[1285] = 8'h81;
Memory[1284] = 8'hB3;
Memory[1291] = 8'h08;
Memory[1290] = 8'h3B;
Memory[1289] = 8'h2C;
Memory[1288] = 8'h23;
Memory[1295] = 8'h00;
Memory[1294] = 8'h80;
Memory[1293] = 8'h01;
Memory[1292] = 8'h13;
Memory[1299] = 8'h00;
Memory[1298] = 8'h0E;
Memory[1297] = 8'h8E;
Memory[1296] = 8'h13;
Memory[1303] = 8'h18;
Memory[1302] = 8'h00;
Memory[1301] = 8'h0A;
Memory[1300] = 8'h63;
Memory[1307] = 8'h00;
Memory[1306] = 8'h50;
Memory[1305] = 8'h01;
Memory[1304] = 8'h13;
Memory[1311] = 8'h0C;
Memory[1310] = 8'h8B;
Memory[1309] = 8'h21;
Memory[1308] = 8'h83;
Memory[1315] = 8'h0C;
Memory[1314] = 8'hCB;
Memory[1313] = 8'h22;
Memory[1312] = 8'h03;
Memory[1319] = 8'h00;
Memory[1318] = 8'h3B;
Memory[1317] = 8'h20;
Memory[1316] = 8'h23;
Memory[1323] = 8'h00;
Memory[1322] = 8'h4B;
Memory[1321] = 8'h22;
Memory[1320] = 8'h23;
Memory[1327] = 8'h01;
Memory[1326] = 8'hDE;
Memory[1325] = 8'h14;
Memory[1324] = 8'h63;
Memory[1331] = 8'h09;
Memory[1330] = 8'hC0;
Memory[1329] = 8'h00;
Memory[1328] = 8'h6F;
Memory[1335] = 8'h01;
Memory[1334] = 8'hDE;
Memory[1333] = 8'h42;
Memory[1332] = 8'h33;
Memory[1339] = 8'h01;
Memory[1338] = 8'h82;
Memory[1337] = 8'h71;
Memory[1336] = 8'hB3;
Memory[1343] = 8'h01;
Memory[1342] = 8'hD1;
Memory[1341] = 8'hF1;
Memory[1340] = 8'hB3;
Memory[1347] = 8'h00;
Memory[1346] = 8'h01;
Memory[1345] = 8'h84;
Memory[1344] = 8'h63;
Memory[1351] = 8'h0D;
Memory[1350] = 8'h00;
Memory[1349] = 8'h21;
Memory[1348] = 8'hEF;
Memory[1355] = 8'hFF;
Memory[1354] = 8'hF2;
Memory[1353] = 8'h71;
Memory[1352] = 8'h93;
Memory[1359] = 8'h01;
Memory[1358] = 8'hD1;
Memory[1357] = 8'hF1;
Memory[1356] = 8'hB3;
Memory[1363] = 8'hD6;
Memory[1362] = 8'h01;
Memory[1361] = 8'h8A;
Memory[1360] = 8'hE3;
Memory[1367] = 8'h40;
Memory[1366] = 8'h01;
Memory[1365] = 8'hF2;
Memory[1364] = 8'h13;
Memory[1371] = 8'h00;
Memory[1370] = 8'h02;
Memory[1369] = 8'h1C;
Memory[1368] = 8'h63;
Memory[1375] = 8'h01;
Memory[1374] = 8'h01;
Memory[1373] = 8'hF2;
Memory[1372] = 8'h13;
Memory[1379] = 8'h00;
Memory[1378] = 8'h02;
Memory[1377] = 8'h1E;
Memory[1376] = 8'h63;
Memory[1383] = 8'h00;
Memory[1382] = 8'h41;
Memory[1381] = 8'hF2;
Memory[1380] = 8'h13;
Memory[1387] = 8'h02;
Memory[1386] = 8'h02;
Memory[1385] = 8'h10;
Memory[1384] = 8'h63;
Memory[1391] = 8'h2C;
Memory[1390] = 8'h40;
Memory[1389] = 8'h00;
Memory[1388] = 8'h6F;
Memory[1395] = 8'h00;
Memory[1394] = 8'h40;
Memory[1393] = 8'h01;
Memory[1392] = 8'h13;
Memory[1399] = 8'h00;
Memory[1398] = 8'h0E;
Memory[1397] = 8'h8E;
Memory[1396] = 8'h13;
Memory[1403] = 8'hF0;
Memory[1402] = 8'h00;
Memory[1401] = 8'h0A;
Memory[1400] = 8'hE3;
Memory[1407] = 8'h00;
Memory[1406] = 8'h60;
Memory[1405] = 8'h01;
Memory[1404] = 8'h13;
Memory[1411] = 8'h00;
Memory[1410] = 8'h0E;
Memory[1409] = 8'h8E;
Memory[1408] = 8'h13;
Memory[1415] = 8'h02;
Memory[1414] = 8'h00;
Memory[1413] = 8'h00;
Memory[1412] = 8'h63;
Memory[1419] = 8'h06;
Memory[1418] = 8'h40;
Memory[1417] = 8'h01;
Memory[1416] = 8'h93;
Memory[1423] = 8'h03;
Memory[1422] = 8'hB1;
Memory[1421] = 8'h81;
Memory[1420] = 8'hB3;
Memory[1427] = 8'h03;
Memory[1426] = 8'hB1;
Memory[1425] = 8'h81;
Memory[1424] = 8'hB3;
Memory[1431] = 8'h08;
Memory[1430] = 8'h3B;
Memory[1429] = 8'h2C;
Memory[1428] = 8'h23;
Memory[1435] = 8'h00;
Memory[1434] = 8'h80;
Memory[1433] = 8'h01;
Memory[1432] = 8'h13;
Memory[1439] = 8'h00;
Memory[1438] = 8'h0E;
Memory[1437] = 8'h8E;
Memory[1436] = 8'h13;
Memory[1443] = 8'h10;
Memory[1442] = 8'h00;
Memory[1441] = 8'h04;
Memory[1440] = 8'h63;
Memory[1447] = 8'h00;
Memory[1446] = 8'h60;
Memory[1445] = 8'h01;
Memory[1444] = 8'h13;
Memory[1451] = 8'h0D;
Memory[1450] = 8'h0B;
Memory[1449] = 8'h21;
Memory[1448] = 8'h83;
Memory[1455] = 8'h0D;
Memory[1454] = 8'h4B;
Memory[1453] = 8'h22;
Memory[1452] = 8'h03;
Memory[1459] = 8'h00;
Memory[1458] = 8'h3B;
Memory[1457] = 8'h20;
Memory[1456] = 8'h23;
Memory[1463] = 8'h00;
Memory[1462] = 8'h4B;
Memory[1461] = 8'h22;
Memory[1460] = 8'h23;
Memory[1467] = 8'h01;
Memory[1466] = 8'hDE;
Memory[1465] = 8'h14;
Memory[1464] = 8'h63;
Memory[1471] = 8'h09;
Memory[1470] = 8'hC0;
Memory[1469] = 8'h00;
Memory[1468] = 8'h6F;
Memory[1475] = 8'h01;
Memory[1474] = 8'hDE;
Memory[1473] = 8'h42;
Memory[1472] = 8'h33;
Memory[1479] = 8'h01;
Memory[1478] = 8'h82;
Memory[1477] = 8'h71;
Memory[1476] = 8'hB3;
Memory[1483] = 8'h01;
Memory[1482] = 8'hD1;
Memory[1481] = 8'hF1;
Memory[1480] = 8'hB3;
Memory[1487] = 8'h00;
Memory[1486] = 8'h01;
Memory[1485] = 8'h84;
Memory[1484] = 8'h63;
Memory[1491] = 8'h0D;
Memory[1490] = 8'h00;
Memory[1489] = 8'h20;
Memory[1488] = 8'h6F;
Memory[1495] = 8'hFF;
Memory[1494] = 8'hF2;
Memory[1493] = 8'h71;
Memory[1492] = 8'h93;
Memory[1499] = 8'h01;
Memory[1498] = 8'hD1;
Memory[1497] = 8'hF1;
Memory[1496] = 8'hB3;
Memory[1503] = 8'hCE;
Memory[1502] = 8'h01;
Memory[1501] = 8'h84;
Memory[1500] = 8'hE3;
Memory[1507] = 8'h40;
Memory[1506] = 8'h01;
Memory[1505] = 8'hF2;
Memory[1504] = 8'h13;
Memory[1511] = 8'hF0;
Memory[1510] = 8'h02;
Memory[1509] = 8'h10;
Memory[1508] = 8'hE3;
Memory[1515] = 8'h01;
Memory[1514] = 8'h01;
Memory[1513] = 8'hF2;
Memory[1512] = 8'h13;
Memory[1519] = 8'hF0;
Memory[1518] = 8'h02;
Memory[1517] = 8'h12;
Memory[1516] = 8'hE3;
Memory[1523] = 8'h00;
Memory[1522] = 8'h41;
Memory[1521] = 8'hF2;
Memory[1520] = 8'h13;
Memory[1527] = 8'hF0;
Memory[1526] = 8'h02;
Memory[1525] = 8'h14;
Memory[1524] = 8'hE3;
Memory[1531] = 8'h2C;
Memory[1530] = 8'h40;
Memory[1529] = 8'h00;
Memory[1528] = 8'h6F;
Memory[1535] = 8'h00;
Memory[1534] = 8'h50;
Memory[1533] = 8'h01;
Memory[1532] = 8'h13;
Memory[1539] = 8'h00;
Memory[1538] = 8'h0E;
Memory[1537] = 8'h8E;
Memory[1536] = 8'h13;
Memory[1543] = 8'hF0;
Memory[1542] = 8'h00;
Memory[1541] = 8'h0A;
Memory[1540] = 8'hE3;
Memory[1547] = 8'h00;
Memory[1546] = 8'h70;
Memory[1545] = 8'h01;
Memory[1544] = 8'h13;
Memory[1551] = 8'h00;
Memory[1550] = 8'h0E;
Memory[1549] = 8'h8E;
Memory[1548] = 8'h13;
Memory[1555] = 8'h02;
Memory[1554] = 8'h00;
Memory[1553] = 8'h00;
Memory[1552] = 8'h63;
Memory[1559] = 8'h1F;
Memory[1558] = 8'h40;
Memory[1557] = 8'h01;
Memory[1556] = 8'h93;
Memory[1563] = 8'h03;
Memory[1562] = 8'hB1;
Memory[1561] = 8'h81;
Memory[1560] = 8'hB3;
Memory[1567] = 8'h03;
Memory[1566] = 8'hB1;
Memory[1565] = 8'h81;
Memory[1564] = 8'hB3;
Memory[1571] = 8'h08;
Memory[1570] = 8'h3B;
Memory[1569] = 8'h2C;
Memory[1568] = 8'h23;
Memory[1575] = 8'h00;
Memory[1574] = 8'h80;
Memory[1573] = 8'h01;
Memory[1572] = 8'h13;
Memory[1579] = 8'h00;
Memory[1578] = 8'h0E;
Memory[1577] = 8'h8E;
Memory[1576] = 8'h13;
Memory[1583] = 8'h06;
Memory[1582] = 8'h00;
Memory[1581] = 8'h0E;
Memory[1580] = 8'h63;
Memory[1587] = 8'h00;
Memory[1586] = 8'h70;
Memory[1585] = 8'h01;
Memory[1584] = 8'h13;
Memory[1591] = 8'h0D;
Memory[1590] = 8'h8B;
Memory[1589] = 8'h21;
Memory[1588] = 8'h83;
Memory[1595] = 8'h0D;
Memory[1594] = 8'hCB;
Memory[1593] = 8'h22;
Memory[1592] = 8'h03;
Memory[1599] = 8'h00;
Memory[1598] = 8'h3B;
Memory[1597] = 8'h20;
Memory[1596] = 8'h23;
Memory[1603] = 8'h00;
Memory[1602] = 8'h4B;
Memory[1601] = 8'h22;
Memory[1600] = 8'h23;
Memory[1607] = 8'h01;
Memory[1606] = 8'hDE;
Memory[1605] = 8'h14;
Memory[1604] = 8'h63;
Memory[1611] = 8'h09;
Memory[1610] = 8'hC0;
Memory[1609] = 8'h00;
Memory[1608] = 8'h6F;
Memory[1615] = 8'h01;
Memory[1614] = 8'hDE;
Memory[1613] = 8'h42;
Memory[1612] = 8'h33;
Memory[1619] = 8'h01;
Memory[1618] = 8'h82;
Memory[1617] = 8'h71;
Memory[1616] = 8'hB3;
Memory[1623] = 8'h01;
Memory[1622] = 8'hD1;
Memory[1621] = 8'hF1;
Memory[1620] = 8'hB3;
Memory[1627] = 8'h00;
Memory[1626] = 8'h01;
Memory[1625] = 8'h84;
Memory[1624] = 8'h63;
Memory[1631] = 8'h0D;
Memory[1630] = 8'h00;
Memory[1629] = 8'h20;
Memory[1628] = 8'h6F;
Memory[1635] = 8'hFF;
Memory[1634] = 8'hF2;
Memory[1633] = 8'h71;
Memory[1632] = 8'h93;
Memory[1639] = 8'h01;
Memory[1638] = 8'hD1;
Memory[1637] = 8'hF1;
Memory[1636] = 8'hB3;
Memory[1643] = 8'hC4;
Memory[1642] = 8'h01;
Memory[1641] = 8'h8E;
Memory[1640] = 8'hE3;
Memory[1647] = 8'h40;
Memory[1646] = 8'h01;
Memory[1645] = 8'hF2;
Memory[1644] = 8'h13;
Memory[1651] = 8'hE6;
Memory[1650] = 8'h02;
Memory[1649] = 8'h1A;
Memory[1648] = 8'hE3;
Memory[1655] = 8'h00;
Memory[1654] = 8'h41;
Memory[1653] = 8'hF2;
Memory[1652] = 8'h13;
Memory[1659] = 8'hE8;
Memory[1658] = 8'h02;
Memory[1657] = 8'h12;
Memory[1656] = 8'hE3;
Memory[1663] = 8'hC4;
Memory[1662] = 8'h00;
Memory[1661] = 8'h04;
Memory[1660] = 8'hE3;
Memory[1667] = 8'h00;
Memory[1666] = 8'h60;
Memory[1665] = 8'h01;
Memory[1664] = 8'h13;
Memory[1671] = 8'h00;
Memory[1670] = 8'h0E;
Memory[1669] = 8'h8E;
Memory[1668] = 8'h13;
Memory[1675] = 8'hF0;
Memory[1674] = 8'h00;
Memory[1673] = 8'h0E;
Memory[1672] = 8'hE3;
Memory[1679] = 8'h3E;
Memory[1678] = 8'h80;
Memory[1677] = 8'h01;
Memory[1676] = 8'h93;
Memory[1683] = 8'h03;
Memory[1682] = 8'hB1;
Memory[1681] = 8'h81;
Memory[1680] = 8'hB3;
Memory[1687] = 8'h03;
Memory[1686] = 8'hB1;
Memory[1685] = 8'h81;
Memory[1684] = 8'hB3;
Memory[1691] = 8'h08;
Memory[1690] = 8'h3B;
Memory[1689] = 8'h2C;
Memory[1688] = 8'h23;
Memory[1695] = 8'h00;
Memory[1694] = 8'h80;
Memory[1693] = 8'h01;
Memory[1692] = 8'h13;
Memory[1699] = 8'h00;
Memory[1698] = 8'h0E;
Memory[1697] = 8'h8E;
Memory[1696] = 8'h13;
Memory[1703] = 8'h00;
Memory[1702] = 8'h00;
Memory[1701] = 8'h02;
Memory[1700] = 8'h63;
Memory[1707] = 8'h00;
Memory[1706] = 8'h80;
Memory[1705] = 8'h01;
Memory[1704] = 8'h13;
Memory[1711] = 8'h0E;
Memory[1710] = 8'h0B;
Memory[1709] = 8'h21;
Memory[1708] = 8'h83;
Memory[1715] = 8'h0E;
Memory[1714] = 8'h4B;
Memory[1713] = 8'h22;
Memory[1712] = 8'h03;
Memory[1719] = 8'h01;
Memory[1718] = 8'hB0;
Memory[1717] = 8'h02;
Memory[1716] = 8'h93;
Memory[1723] = 8'h00;
Memory[1722] = 8'h3B;
Memory[1721] = 8'h20;
Memory[1720] = 8'h23;
Memory[1727] = 8'h00;
Memory[1726] = 8'h4B;
Memory[1725] = 8'h22;
Memory[1724] = 8'h23;
Memory[1731] = 8'h00;
Memory[1730] = 8'h5B;
Memory[1729] = 8'h24;
Memory[1728] = 8'h23;
Memory[1735] = 8'h01;
Memory[1734] = 8'hDE;
Memory[1733] = 8'h14;
Memory[1732] = 8'h63;
Memory[1739] = 8'h09;
Memory[1738] = 8'hC0;
Memory[1737] = 8'h00;
Memory[1736] = 8'h6F;
Memory[1743] = 8'h01;
Memory[1742] = 8'hDE;
Memory[1741] = 8'h42;
Memory[1740] = 8'h33;
Memory[1747] = 8'h01;
Memory[1746] = 8'h82;
Memory[1745] = 8'h71;
Memory[1744] = 8'hB3;
Memory[1751] = 8'h01;
Memory[1750] = 8'hD1;
Memory[1749] = 8'hF1;
Memory[1748] = 8'hB3;
Memory[1755] = 8'h00;
Memory[1754] = 8'h01;
Memory[1753] = 8'h84;
Memory[1752] = 8'h63;
Memory[1759] = 8'h0D;
Memory[1758] = 8'h00;
Memory[1757] = 8'h20;
Memory[1756] = 8'h6F;
Memory[1763] = 8'hFF;
Memory[1762] = 8'hF2;
Memory[1761] = 8'h71;
Memory[1760] = 8'h93;
Memory[1767] = 8'h01;
Memory[1766] = 8'hD1;
Memory[1765] = 8'hF1;
Memory[1764] = 8'hB3;
Memory[1771] = 8'hBC;
Memory[1770] = 8'h01;
Memory[1769] = 8'h8E;
Memory[1768] = 8'hE3;
Memory[1775] = 8'h04;
Memory[1774] = 8'h01;
Memory[1773] = 8'hF2;
Memory[1772] = 8'h13;
Memory[1779] = 8'h00;
Memory[1778] = 8'h02;
Memory[1777] = 8'h18;
Memory[1776] = 8'h63;
Memory[1783] = 8'h00;
Memory[1782] = 8'h41;
Memory[1781] = 8'hF2;
Memory[1780] = 8'h13;
Memory[1787] = 8'h00;
Memory[1786] = 8'h02;
Memory[1785] = 8'h1A;
Memory[1784] = 8'h63;
Memory[1791] = 8'h2C;
Memory[1790] = 8'h40;
Memory[1789] = 8'h00;
Memory[1788] = 8'h6F;
Memory[1795] = 8'h00;
Memory[1794] = 8'h90;
Memory[1793] = 8'h01;
Memory[1792] = 8'h13;
Memory[1799] = 8'h00;
Memory[1798] = 8'h0E;
Memory[1797] = 8'h8E;
Memory[1796] = 8'h13;
Memory[1803] = 8'h00;
Memory[1802] = 8'h00;
Memory[1801] = 8'h08;
Memory[1800] = 8'h63;
Memory[1807] = 8'h02;
Memory[1806] = 8'h50;
Memory[1805] = 8'h01;
Memory[1804] = 8'h13;
Memory[1811] = 8'h00;
Memory[1810] = 8'h0E;
Memory[1809] = 8'h8E;
Memory[1808] = 8'h13;
Memory[1815] = 8'h67;
Memory[1814] = 8'h40;
Memory[1813] = 8'h10;
Memory[1812] = 8'h6F;
Memory[1819] = 8'h00;
Memory[1818] = 8'h90;
Memory[1817] = 8'h01;
Memory[1816] = 8'h13;
Memory[1823] = 8'h0E;
Memory[1822] = 8'h8B;
Memory[1821] = 8'h21;
Memory[1820] = 8'h83;
Memory[1827] = 8'h0E;
Memory[1826] = 8'hCB;
Memory[1825] = 8'h22;
Memory[1824] = 8'h03;
Memory[1831] = 8'h01;
Memory[1830] = 8'hB0;
Memory[1829] = 8'h02;
Memory[1828] = 8'h93;
Memory[1835] = 8'h00;
Memory[1834] = 8'h3B;
Memory[1833] = 8'h20;
Memory[1832] = 8'h23;
Memory[1839] = 8'h00;
Memory[1838] = 8'h4B;
Memory[1837] = 8'h22;
Memory[1836] = 8'h23;
Memory[1843] = 8'h00;
Memory[1842] = 8'h5B;
Memory[1841] = 8'h24;
Memory[1840] = 8'h23;
Memory[1847] = 8'h01;
Memory[1846] = 8'hDE;
Memory[1845] = 8'h14;
Memory[1844] = 8'h63;
Memory[1851] = 8'h09;
Memory[1850] = 8'hC0;
Memory[1849] = 8'h00;
Memory[1848] = 8'h6F;
Memory[1855] = 8'h01;
Memory[1854] = 8'hDE;
Memory[1853] = 8'h42;
Memory[1852] = 8'h33;
Memory[1859] = 8'h01;
Memory[1858] = 8'h82;
Memory[1857] = 8'h71;
Memory[1856] = 8'hB3;
Memory[1863] = 8'h01;
Memory[1862] = 8'hD1;
Memory[1861] = 8'hF1;
Memory[1860] = 8'hB3;
Memory[1867] = 8'h00;
Memory[1866] = 8'h01;
Memory[1865] = 8'h84;
Memory[1864] = 8'h63;
Memory[1871] = 8'h0D;
Memory[1870] = 8'h00;
Memory[1869] = 8'h20;
Memory[1868] = 8'h6F;
Memory[1875] = 8'hFF;
Memory[1874] = 8'hF2;
Memory[1873] = 8'h71;
Memory[1872] = 8'h93;
Memory[1879] = 8'h01;
Memory[1878] = 8'hD1;
Memory[1877] = 8'hF1;
Memory[1876] = 8'hB3;
Memory[1883] = 8'hB6;
Memory[1882] = 8'h01;
Memory[1881] = 8'h86;
Memory[1880] = 8'hE3;
Memory[1887] = 8'h10;
Memory[1886] = 8'h01;
Memory[1885] = 8'hF2;
Memory[1884] = 8'h13;
Memory[1891] = 8'h00;
Memory[1890] = 8'h02;
Memory[1889] = 8'h1C;
Memory[1888] = 8'h63;
Memory[1895] = 8'h04;
Memory[1894] = 8'h01;
Memory[1893] = 8'hF2;
Memory[1892] = 8'h13;
Memory[1899] = 8'h00;
Memory[1898] = 8'h02;
Memory[1897] = 8'h1E;
Memory[1896] = 8'h63;
Memory[1903] = 8'h00;
Memory[1902] = 8'h41;
Memory[1901] = 8'hF2;
Memory[1900] = 8'h13;
Memory[1907] = 8'h02;
Memory[1906] = 8'h02;
Memory[1905] = 8'h10;
Memory[1904] = 8'h63;
Memory[1911] = 8'hB4;
Memory[1910] = 8'h00;
Memory[1909] = 8'h08;
Memory[1908] = 8'hE3;
Memory[1915] = 8'h00;
Memory[1914] = 8'h80;
Memory[1913] = 8'h01;
Memory[1912] = 8'h13;
Memory[1919] = 8'h00;
Memory[1918] = 8'h0E;
Memory[1917] = 8'h8E;
Memory[1916] = 8'h13;
Memory[1923] = 8'hF2;
Memory[1922] = 8'h00;
Memory[1921] = 8'h04;
Memory[1920] = 8'hE3;
Memory[1927] = 8'h01;
Memory[1926] = 8'h30;
Memory[1925] = 8'h01;
Memory[1924] = 8'h13;
Memory[1931] = 8'h00;
Memory[1930] = 8'h0E;
Memory[1929] = 8'h8E;
Memory[1928] = 8'h13;
Memory[1935] = 8'h3E;
Memory[1934] = 8'h00;
Memory[1933] = 8'h04;
Memory[1932] = 8'h63;
Memory[1939] = 8'h00;
Memory[1938] = 8'hA0;
Memory[1937] = 8'h01;
Memory[1936] = 8'h13;
Memory[1943] = 8'h00;
Memory[1942] = 8'h0E;
Memory[1941] = 8'h8E;
Memory[1940] = 8'h13;
Memory[1947] = 8'h00;
Memory[1946] = 8'h00;
Memory[1945] = 8'h02;
Memory[1944] = 8'h63;
Memory[1951] = 8'h00;
Memory[1950] = 8'hA0;
Memory[1949] = 8'h01;
Memory[1948] = 8'h13;
Memory[1955] = 8'h0F;
Memory[1954] = 8'h0B;
Memory[1953] = 8'h21;
Memory[1952] = 8'h83;
Memory[1959] = 8'h07;
Memory[1958] = 8'h4B;
Memory[1957] = 8'h23;
Memory[1956] = 8'h83;
Memory[1963] = 8'h06;
Memory[1962] = 8'h40;
Memory[1961] = 8'h02;
Memory[1960] = 8'h93;
Memory[1967] = 8'h03;
Memory[1966] = 8'hB2;
Memory[1965] = 8'h82;
Memory[1964] = 8'hB3;
Memory[1971] = 8'h02;
Memory[1970] = 8'h53;
Memory[1969] = 8'hC2;
Memory[1968] = 8'h33;
Memory[1975] = 8'h00;
Memory[1974] = 8'hA0;
Memory[1973] = 8'h02;
Memory[1972] = 8'h93;
Memory[1979] = 8'h02;
Memory[1978] = 8'h52;
Memory[1977] = 8'h62;
Memory[1976] = 8'h33;
Memory[1983] = 8'h00;
Memory[1982] = 8'h82;
Memory[1981] = 8'h12;
Memory[1980] = 8'h13;
Memory[1987] = 8'h00;
Memory[1986] = 8'hA0;
Memory[1985] = 8'h02;
Memory[1984] = 8'h93;
Memory[1991] = 8'h03;
Memory[1990] = 8'hB2;
Memory[1989] = 8'h82;
Memory[1988] = 8'hB3;
Memory[1995] = 8'h02;
Memory[1994] = 8'h53;
Memory[1993] = 8'hC3;
Memory[1992] = 8'h33;
Memory[1999] = 8'h00;
Memory[1998] = 8'hA0;
Memory[1997] = 8'h02;
Memory[1996] = 8'h93;
Memory[2003] = 8'h02;
Memory[2002] = 8'h53;
Memory[2001] = 8'h63;
Memory[2000] = 8'h33;
Memory[2007] = 8'h00;
Memory[2006] = 8'h62;
Memory[2005] = 8'h02;
Memory[2004] = 8'h33;
Memory[2011] = 8'h00;
Memory[2010] = 8'h41;
Memory[2009] = 8'h81;
Memory[2008] = 8'hB3;
Memory[2015] = 8'h00;
Memory[2014] = 8'h3B;
Memory[2013] = 8'h20;
Memory[2012] = 8'h23;
Memory[2019] = 8'h0F;
Memory[2018] = 8'h4B;
Memory[2017] = 8'h21;
Memory[2016] = 8'h83;
Memory[2023] = 8'h3E;
Memory[2022] = 8'h80;
Memory[2021] = 8'h02;
Memory[2020] = 8'h93;
Memory[2027] = 8'h02;
Memory[2026] = 8'h53;
Memory[2025] = 8'hC2;
Memory[2024] = 8'h33;
Memory[2031] = 8'h00;
Memory[2030] = 8'hA0;
Memory[2029] = 8'h02;
Memory[2028] = 8'h93;
Memory[2035] = 8'h02;
Memory[2034] = 8'h52;
Memory[2033] = 8'h62;
Memory[2032] = 8'h33;
Memory[2039] = 8'h00;
Memory[2038] = 8'h82;
Memory[2037] = 8'h12;
Memory[2036] = 8'h13;
Memory[2043] = 8'h06;
Memory[2042] = 8'h40;
Memory[2041] = 8'h02;
Memory[2040] = 8'h93;
Memory[2047] = 8'h02;
Memory[2046] = 8'h53;
Memory[2045] = 8'hC3;
Memory[2044] = 8'h33;
Memory[2051] = 8'h00;
Memory[2050] = 8'hA0;
Memory[2049] = 8'h02;
Memory[2048] = 8'h93;
Memory[2055] = 8'h02;
Memory[2054] = 8'h53;
Memory[2053] = 8'h63;
Memory[2052] = 8'h33;
Memory[2059] = 8'h00;
Memory[2058] = 8'h62;
Memory[2057] = 8'h02;
Memory[2056] = 8'h33;
Memory[2063] = 8'h00;
Memory[2062] = 8'h82;
Memory[2061] = 8'h12;
Memory[2060] = 8'h13;
Memory[2067] = 8'h02;
Memory[2066] = 8'h53;
Memory[2065] = 8'hC3;
Memory[2064] = 8'h33;
Memory[2071] = 8'h02;
Memory[2070] = 8'h53;
Memory[2069] = 8'h63;
Memory[2068] = 8'h33;
Memory[2075] = 8'h00;
Memory[2074] = 8'h62;
Memory[2073] = 8'h02;
Memory[2072] = 8'h33;
Memory[2079] = 8'h00;
Memory[2078] = 8'h82;
Memory[2077] = 8'h12;
Memory[2076] = 8'h13;
Memory[2083] = 8'h02;
Memory[2082] = 8'h53;
Memory[2081] = 8'hE3;
Memory[2080] = 8'h33;
Memory[2087] = 8'h00;
Memory[2086] = 8'h62;
Memory[2085] = 8'h02;
Memory[2084] = 8'h33;
Memory[2091] = 8'h00;
Memory[2090] = 8'h41;
Memory[2089] = 8'h81;
Memory[2088] = 8'hB3;
Memory[2095] = 8'h00;
Memory[2094] = 8'h3B;
Memory[2093] = 8'h22;
Memory[2092] = 8'h23;
Memory[2099] = 8'h01;
Memory[2098] = 8'hDE;
Memory[2097] = 8'h14;
Memory[2096] = 8'h63;
Memory[2103] = 8'h09;
Memory[2102] = 8'hC0;
Memory[2101] = 8'h00;
Memory[2100] = 8'h6F;
Memory[2107] = 8'h01;
Memory[2106] = 8'hDE;
Memory[2105] = 8'h42;
Memory[2104] = 8'h33;
Memory[2111] = 8'h01;
Memory[2110] = 8'h82;
Memory[2109] = 8'h71;
Memory[2108] = 8'hB3;
Memory[2115] = 8'h01;
Memory[2114] = 8'hD1;
Memory[2113] = 8'hF1;
Memory[2112] = 8'hB3;
Memory[2119] = 8'h00;
Memory[2118] = 8'h01;
Memory[2117] = 8'h84;
Memory[2116] = 8'h63;
Memory[2123] = 8'h0D;
Memory[2122] = 8'h00;
Memory[2121] = 8'h20;
Memory[2120] = 8'h6F;
Memory[2127] = 8'hFF;
Memory[2126] = 8'hF2;
Memory[2125] = 8'h71;
Memory[2124] = 8'h93;
Memory[2131] = 8'h01;
Memory[2130] = 8'hD1;
Memory[2129] = 8'hF1;
Memory[2128] = 8'hB3;
Memory[2135] = 8'h00;
Memory[2134] = 8'h01;
Memory[2133] = 8'h94;
Memory[2132] = 8'h63;
Memory[2139] = 8'h2C;
Memory[2138] = 8'h40;
Memory[2137] = 8'h00;
Memory[2136] = 8'h6F;
Memory[2143] = 8'h04;
Memory[2142] = 8'h01;
Memory[2141] = 8'hF2;
Memory[2140] = 8'h13;
Memory[2147] = 8'h00;
Memory[2146] = 8'h02;
Memory[2145] = 8'h18;
Memory[2144] = 8'h63;
Memory[2151] = 8'h00;
Memory[2150] = 8'h11;
Memory[2149] = 8'hF2;
Memory[2148] = 8'h13;
Memory[2155] = 8'h00;
Memory[2154] = 8'h02;
Memory[2153] = 8'h1A;
Memory[2152] = 8'h63;
Memory[2159] = 8'h2C;
Memory[2158] = 8'h40;
Memory[2157] = 8'h00;
Memory[2156] = 8'h6F;
Memory[2163] = 8'h00;
Memory[2162] = 8'hB0;
Memory[2161] = 8'h01;
Memory[2160] = 8'h13;
Memory[2167] = 8'h00;
Memory[2166] = 8'h0E;
Memory[2165] = 8'h8E;
Memory[2164] = 8'h13;
Memory[2171] = 8'h08;
Memory[2170] = 8'h90;
Memory[2169] = 8'h00;
Memory[2168] = 8'h6F;
Memory[2175] = 8'h00;
Memory[2174] = 8'h90;
Memory[2173] = 8'h01;
Memory[2172] = 8'h13;
Memory[2179] = 8'h00;
Memory[2178] = 8'h0E;
Memory[2177] = 8'h8E;
Memory[2176] = 8'h13;
Memory[2183] = 8'h71;
Memory[2182] = 8'h80;
Memory[2181] = 8'h00;
Memory[2180] = 8'h6F;
Memory[2187] = 8'h00;
Memory[2186] = 8'hB0;
Memory[2185] = 8'h01;
Memory[2184] = 8'h13;
Memory[2191] = 8'h0F;
Memory[2190] = 8'h8B;
Memory[2189] = 8'h21;
Memory[2188] = 8'h83;
Memory[2195] = 8'h07;
Memory[2194] = 8'h8B;
Memory[2193] = 8'h23;
Memory[2192] = 8'h83;
Memory[2199] = 8'h06;
Memory[2198] = 8'h40;
Memory[2197] = 8'h02;
Memory[2196] = 8'h93;
Memory[2203] = 8'h03;
Memory[2202] = 8'hB2;
Memory[2201] = 8'h82;
Memory[2200] = 8'hB3;
Memory[2207] = 8'h02;
Memory[2206] = 8'h53;
Memory[2205] = 8'hC2;
Memory[2204] = 8'h33;
Memory[2211] = 8'h00;
Memory[2210] = 8'hA0;
Memory[2209] = 8'h02;
Memory[2208] = 8'h93;
Memory[2215] = 8'h02;
Memory[2214] = 8'h52;
Memory[2213] = 8'h62;
Memory[2212] = 8'h33;
Memory[2219] = 8'h00;
Memory[2218] = 8'h82;
Memory[2217] = 8'h12;
Memory[2216] = 8'h13;
Memory[2223] = 8'h00;
Memory[2222] = 8'hA0;
Memory[2221] = 8'h02;
Memory[2220] = 8'h93;
Memory[2227] = 8'h03;
Memory[2226] = 8'hB2;
Memory[2225] = 8'h82;
Memory[2224] = 8'hB3;
Memory[2231] = 8'h02;
Memory[2230] = 8'h53;
Memory[2229] = 8'hC3;
Memory[2228] = 8'h33;
Memory[2235] = 8'h00;
Memory[2234] = 8'hA0;
Memory[2233] = 8'h02;
Memory[2232] = 8'h93;
Memory[2239] = 8'h02;
Memory[2238] = 8'h53;
Memory[2237] = 8'h63;
Memory[2236] = 8'h33;
Memory[2243] = 8'h00;
Memory[2242] = 8'h62;
Memory[2241] = 8'h02;
Memory[2240] = 8'h33;
Memory[2247] = 8'h00;
Memory[2246] = 8'h41;
Memory[2245] = 8'h81;
Memory[2244] = 8'hB3;
Memory[2251] = 8'h00;
Memory[2250] = 8'h3B;
Memory[2249] = 8'h20;
Memory[2248] = 8'h23;
Memory[2255] = 8'h0F;
Memory[2254] = 8'hCB;
Memory[2253] = 8'h21;
Memory[2252] = 8'h83;
Memory[2259] = 8'h3E;
Memory[2258] = 8'h80;
Memory[2257] = 8'h02;
Memory[2256] = 8'h93;
Memory[2263] = 8'h02;
Memory[2262] = 8'h53;
Memory[2261] = 8'hC2;
Memory[2260] = 8'h33;
Memory[2267] = 8'h00;
Memory[2266] = 8'hA0;
Memory[2265] = 8'h02;
Memory[2264] = 8'h93;
Memory[2271] = 8'h02;
Memory[2270] = 8'h52;
Memory[2269] = 8'h62;
Memory[2268] = 8'h33;
Memory[2275] = 8'h00;
Memory[2274] = 8'h82;
Memory[2273] = 8'h12;
Memory[2272] = 8'h13;
Memory[2279] = 8'h06;
Memory[2278] = 8'h40;
Memory[2277] = 8'h02;
Memory[2276] = 8'h93;
Memory[2283] = 8'h02;
Memory[2282] = 8'h53;
Memory[2281] = 8'hC3;
Memory[2280] = 8'h33;
Memory[2287] = 8'h00;
Memory[2286] = 8'hA0;
Memory[2285] = 8'h02;
Memory[2284] = 8'h93;
Memory[2291] = 8'h02;
Memory[2290] = 8'h53;
Memory[2289] = 8'h63;
Memory[2288] = 8'h33;
Memory[2295] = 8'h00;
Memory[2294] = 8'h62;
Memory[2293] = 8'h02;
Memory[2292] = 8'h33;
Memory[2299] = 8'h00;
Memory[2298] = 8'h82;
Memory[2297] = 8'h12;
Memory[2296] = 8'h13;
Memory[2303] = 8'h02;
Memory[2302] = 8'h53;
Memory[2301] = 8'hC3;
Memory[2300] = 8'h33;
Memory[2307] = 8'h02;
Memory[2306] = 8'h53;
Memory[2305] = 8'h63;
Memory[2304] = 8'h33;
Memory[2311] = 8'h00;
Memory[2310] = 8'h62;
Memory[2309] = 8'h02;
Memory[2308] = 8'h33;
Memory[2315] = 8'h00;
Memory[2314] = 8'h82;
Memory[2313] = 8'h12;
Memory[2312] = 8'h13;
Memory[2319] = 8'h02;
Memory[2318] = 8'h53;
Memory[2317] = 8'hE3;
Memory[2316] = 8'h33;
Memory[2323] = 8'h00;
Memory[2322] = 8'h62;
Memory[2321] = 8'h02;
Memory[2320] = 8'h33;
Memory[2327] = 8'h00;
Memory[2326] = 8'h41;
Memory[2325] = 8'h81;
Memory[2324] = 8'hB3;
Memory[2331] = 8'h00;
Memory[2330] = 8'h3B;
Memory[2329] = 8'h22;
Memory[2328] = 8'h23;
Memory[2335] = 8'h01;
Memory[2334] = 8'hDE;
Memory[2333] = 8'h14;
Memory[2332] = 8'h63;
Memory[2339] = 8'h09;
Memory[2338] = 8'hC0;
Memory[2337] = 8'h00;
Memory[2336] = 8'h6F;
Memory[2343] = 8'h01;
Memory[2342] = 8'hDE;
Memory[2341] = 8'h42;
Memory[2340] = 8'h33;
Memory[2347] = 8'h01;
Memory[2346] = 8'h82;
Memory[2345] = 8'h71;
Memory[2344] = 8'hB3;
Memory[2351] = 8'h01;
Memory[2350] = 8'hD1;
Memory[2349] = 8'hF1;
Memory[2348] = 8'hB3;
Memory[2355] = 8'h00;
Memory[2354] = 8'h01;
Memory[2353] = 8'h84;
Memory[2352] = 8'h63;
Memory[2359] = 8'h0D;
Memory[2358] = 8'h00;
Memory[2357] = 8'h20;
Memory[2356] = 8'h6F;
Memory[2363] = 8'hFF;
Memory[2362] = 8'hF2;
Memory[2361] = 8'h71;
Memory[2360] = 8'h93;
Memory[2367] = 8'h01;
Memory[2366] = 8'hD1;
Memory[2365] = 8'hF1;
Memory[2364] = 8'hB3;
Memory[2371] = 8'h00;
Memory[2370] = 8'h01;
Memory[2369] = 8'h94;
Memory[2368] = 8'h63;
Memory[2375] = 8'h2C;
Memory[2374] = 8'h40;
Memory[2373] = 8'h00;
Memory[2372] = 8'h6F;
Memory[2379] = 8'h10;
Memory[2378] = 8'h01;
Memory[2377] = 8'hF2;
Memory[2376] = 8'h13;
Memory[2383] = 8'h00;
Memory[2382] = 8'h02;
Memory[2381] = 8'h1C;
Memory[2380] = 8'h63;
Memory[2387] = 8'h04;
Memory[2386] = 8'h01;
Memory[2385] = 8'hF2;
Memory[2384] = 8'h13;
Memory[2391] = 8'h00;
Memory[2390] = 8'h02;
Memory[2389] = 8'h1E;
Memory[2388] = 8'h63;
Memory[2395] = 8'h00;
Memory[2394] = 8'h11;
Memory[2393] = 8'hF2;
Memory[2392] = 8'h13;
Memory[2399] = 8'h02;
Memory[2398] = 8'h02;
Memory[2397] = 8'h10;
Memory[2396] = 8'h63;
Memory[2403] = 8'h2C;
Memory[2402] = 8'h40;
Memory[2401] = 8'h00;
Memory[2400] = 8'h6F;
Memory[2407] = 8'h00;
Memory[2406] = 8'hA0;
Memory[2405] = 8'h01;
Memory[2404] = 8'h13;
Memory[2411] = 8'h00;
Memory[2410] = 8'h0E;
Memory[2409] = 8'h8E;
Memory[2408] = 8'h13;
Memory[2415] = 8'h79;
Memory[2414] = 8'hC0;
Memory[2413] = 8'h00;
Memory[2412] = 8'h6F;
Memory[2419] = 8'h00;
Memory[2418] = 8'hC0;
Memory[2417] = 8'h01;
Memory[2416] = 8'h13;
Memory[2423] = 8'h00;
Memory[2422] = 8'h0E;
Memory[2421] = 8'h8E;
Memory[2420] = 8'h13;
Memory[2427] = 8'h18;
Memory[2426] = 8'h90;
Memory[2425] = 8'h00;
Memory[2424] = 8'h6F;
Memory[2431] = 8'h00;
Memory[2430] = 8'h90;
Memory[2429] = 8'h01;
Memory[2428] = 8'h13;
Memory[2435] = 8'h00;
Memory[2434] = 8'h0E;
Memory[2433] = 8'h8E;
Memory[2432] = 8'h13;
Memory[2439] = 8'h71;
Memory[2438] = 8'h80;
Memory[2437] = 8'h00;
Memory[2436] = 8'h6F;
Memory[2443] = 8'h00;
Memory[2442] = 8'hC0;
Memory[2441] = 8'h01;
Memory[2440] = 8'h13;
Memory[2447] = 8'h10;
Memory[2446] = 8'h0B;
Memory[2445] = 8'h21;
Memory[2444] = 8'h83;
Memory[2451] = 8'h07;
Memory[2450] = 8'hCB;
Memory[2449] = 8'h23;
Memory[2448] = 8'h83;
Memory[2455] = 8'h06;
Memory[2454] = 8'h40;
Memory[2453] = 8'h02;
Memory[2452] = 8'h93;
Memory[2459] = 8'h03;
Memory[2458] = 8'hB2;
Memory[2457] = 8'h82;
Memory[2456] = 8'hB3;
Memory[2463] = 8'h02;
Memory[2462] = 8'h53;
Memory[2461] = 8'hC2;
Memory[2460] = 8'h33;
Memory[2467] = 8'h00;
Memory[2466] = 8'hA0;
Memory[2465] = 8'h02;
Memory[2464] = 8'h93;
Memory[2471] = 8'h02;
Memory[2470] = 8'h52;
Memory[2469] = 8'h62;
Memory[2468] = 8'h33;
Memory[2475] = 8'h00;
Memory[2474] = 8'h82;
Memory[2473] = 8'h12;
Memory[2472] = 8'h13;
Memory[2479] = 8'h00;
Memory[2478] = 8'hA0;
Memory[2477] = 8'h02;
Memory[2476] = 8'h93;
Memory[2483] = 8'h03;
Memory[2482] = 8'hB2;
Memory[2481] = 8'h82;
Memory[2480] = 8'hB3;
Memory[2487] = 8'h02;
Memory[2486] = 8'h53;
Memory[2485] = 8'hC3;
Memory[2484] = 8'h33;
Memory[2491] = 8'h00;
Memory[2490] = 8'hA0;
Memory[2489] = 8'h02;
Memory[2488] = 8'h93;
Memory[2495] = 8'h02;
Memory[2494] = 8'h53;
Memory[2493] = 8'h63;
Memory[2492] = 8'h33;
Memory[2499] = 8'h00;
Memory[2498] = 8'h62;
Memory[2497] = 8'h02;
Memory[2496] = 8'h33;
Memory[2503] = 8'h00;
Memory[2502] = 8'h41;
Memory[2501] = 8'h81;
Memory[2500] = 8'hB3;
Memory[2507] = 8'h00;
Memory[2506] = 8'h3B;
Memory[2505] = 8'h20;
Memory[2504] = 8'h23;
Memory[2511] = 8'h10;
Memory[2510] = 8'h4B;
Memory[2509] = 8'h21;
Memory[2508] = 8'h83;
Memory[2515] = 8'h3E;
Memory[2514] = 8'h80;
Memory[2513] = 8'h02;
Memory[2512] = 8'h93;
Memory[2519] = 8'h02;
Memory[2518] = 8'h53;
Memory[2517] = 8'hC2;
Memory[2516] = 8'h33;
Memory[2523] = 8'h00;
Memory[2522] = 8'hA0;
Memory[2521] = 8'h02;
Memory[2520] = 8'h93;
Memory[2527] = 8'h02;
Memory[2526] = 8'h52;
Memory[2525] = 8'h62;
Memory[2524] = 8'h33;
Memory[2531] = 8'h00;
Memory[2530] = 8'h82;
Memory[2529] = 8'h12;
Memory[2528] = 8'h13;
Memory[2535] = 8'h06;
Memory[2534] = 8'h40;
Memory[2533] = 8'h02;
Memory[2532] = 8'h93;
Memory[2539] = 8'h02;
Memory[2538] = 8'h53;
Memory[2537] = 8'hC3;
Memory[2536] = 8'h33;
Memory[2543] = 8'h00;
Memory[2542] = 8'hA0;
Memory[2541] = 8'h02;
Memory[2540] = 8'h93;
Memory[2547] = 8'h02;
Memory[2546] = 8'h53;
Memory[2545] = 8'h63;
Memory[2544] = 8'h33;
Memory[2551] = 8'h00;
Memory[2550] = 8'h62;
Memory[2549] = 8'h02;
Memory[2548] = 8'h33;
Memory[2555] = 8'h00;
Memory[2554] = 8'h82;
Memory[2553] = 8'h12;
Memory[2552] = 8'h13;
Memory[2559] = 8'h02;
Memory[2558] = 8'h53;
Memory[2557] = 8'hC3;
Memory[2556] = 8'h33;
Memory[2563] = 8'h02;
Memory[2562] = 8'h53;
Memory[2561] = 8'h63;
Memory[2560] = 8'h33;
Memory[2567] = 8'h00;
Memory[2566] = 8'h62;
Memory[2565] = 8'h02;
Memory[2564] = 8'h33;
Memory[2571] = 8'h00;
Memory[2570] = 8'h82;
Memory[2569] = 8'h12;
Memory[2568] = 8'h13;
Memory[2575] = 8'h02;
Memory[2574] = 8'h53;
Memory[2573] = 8'hE3;
Memory[2572] = 8'h33;
Memory[2579] = 8'h00;
Memory[2578] = 8'h62;
Memory[2577] = 8'h02;
Memory[2576] = 8'h33;
Memory[2583] = 8'h00;
Memory[2582] = 8'h41;
Memory[2581] = 8'h81;
Memory[2580] = 8'hB3;
Memory[2587] = 8'h00;
Memory[2586] = 8'h3B;
Memory[2585] = 8'h22;
Memory[2584] = 8'h23;
Memory[2591] = 8'h01;
Memory[2590] = 8'hDE;
Memory[2589] = 8'h14;
Memory[2588] = 8'h63;
Memory[2595] = 8'h09;
Memory[2594] = 8'hC0;
Memory[2593] = 8'h00;
Memory[2592] = 8'h6F;
Memory[2599] = 8'h01;
Memory[2598] = 8'hDE;
Memory[2597] = 8'h42;
Memory[2596] = 8'h33;
Memory[2603] = 8'h01;
Memory[2602] = 8'h82;
Memory[2601] = 8'h71;
Memory[2600] = 8'hB3;
Memory[2607] = 8'h01;
Memory[2606] = 8'hD1;
Memory[2605] = 8'hF1;
Memory[2604] = 8'hB3;
Memory[2611] = 8'h00;
Memory[2610] = 8'h01;
Memory[2609] = 8'h84;
Memory[2608] = 8'h63;
Memory[2615] = 8'h0D;
Memory[2614] = 8'h00;
Memory[2613] = 8'h20;
Memory[2612] = 8'h6F;
Memory[2619] = 8'hFF;
Memory[2618] = 8'hF2;
Memory[2617] = 8'h71;
Memory[2616] = 8'h93;
Memory[2623] = 8'h01;
Memory[2622] = 8'hD1;
Memory[2621] = 8'hF1;
Memory[2620] = 8'hB3;
Memory[2627] = 8'h00;
Memory[2626] = 8'h01;
Memory[2625] = 8'h94;
Memory[2624] = 8'h63;
Memory[2631] = 8'h2C;
Memory[2630] = 8'h40;
Memory[2629] = 8'h00;
Memory[2628] = 8'h6F;
Memory[2635] = 8'h10;
Memory[2634] = 8'h01;
Memory[2633] = 8'hF2;
Memory[2632] = 8'h13;
Memory[2639] = 8'h00;
Memory[2638] = 8'h02;
Memory[2637] = 8'h1C;
Memory[2636] = 8'h63;
Memory[2643] = 8'h04;
Memory[2642] = 8'h01;
Memory[2641] = 8'hF2;
Memory[2640] = 8'h13;
Memory[2647] = 8'h00;
Memory[2646] = 8'h02;
Memory[2645] = 8'h1E;
Memory[2644] = 8'h63;
Memory[2651] = 8'h00;
Memory[2650] = 8'h11;
Memory[2649] = 8'hF2;
Memory[2648] = 8'h13;
Memory[2655] = 8'h02;
Memory[2654] = 8'h02;
Memory[2653] = 8'h10;
Memory[2652] = 8'h63;
Memory[2659] = 8'h2C;
Memory[2658] = 8'h40;
Memory[2657] = 8'h00;
Memory[2656] = 8'h6F;
Memory[2663] = 8'h00;
Memory[2662] = 8'hB0;
Memory[2661] = 8'h01;
Memory[2660] = 8'h13;
Memory[2667] = 8'h00;
Memory[2666] = 8'h0E;
Memory[2665] = 8'h8E;
Memory[2664] = 8'h13;
Memory[2671] = 8'h08;
Memory[2670] = 8'h90;
Memory[2669] = 8'h00;
Memory[2668] = 8'h6F;
Memory[2675] = 8'h00;
Memory[2674] = 8'hD0;
Memory[2673] = 8'h01;
Memory[2672] = 8'h13;
Memory[2679] = 8'h00;
Memory[2678] = 8'h0E;
Memory[2677] = 8'h8E;
Memory[2676] = 8'h13;
Memory[2683] = 8'h00;
Memory[2682] = 8'h00;
Memory[2681] = 8'h08;
Memory[2680] = 8'h63;
Memory[2687] = 8'h00;
Memory[2686] = 8'h90;
Memory[2685] = 8'h01;
Memory[2684] = 8'h13;
Memory[2691] = 8'h00;
Memory[2690] = 8'h0E;
Memory[2689] = 8'h8E;
Memory[2688] = 8'h13;
Memory[2695] = 8'h71;
Memory[2694] = 8'h80;
Memory[2693] = 8'h00;
Memory[2692] = 8'h6F;
Memory[2699] = 8'h00;
Memory[2698] = 8'hD0;
Memory[2697] = 8'h01;
Memory[2696] = 8'h13;
Memory[2703] = 8'h10;
Memory[2702] = 8'h8B;
Memory[2701] = 8'h21;
Memory[2700] = 8'h83;
Memory[2707] = 8'h08;
Memory[2706] = 8'h0B;
Memory[2705] = 8'h23;
Memory[2704] = 8'h83;
Memory[2711] = 8'h06;
Memory[2710] = 8'h40;
Memory[2709] = 8'h02;
Memory[2708] = 8'h93;
Memory[2715] = 8'h03;
Memory[2714] = 8'hB2;
Memory[2713] = 8'h82;
Memory[2712] = 8'hB3;
Memory[2719] = 8'h02;
Memory[2718] = 8'h53;
Memory[2717] = 8'hC2;
Memory[2716] = 8'h33;
Memory[2723] = 8'h00;
Memory[2722] = 8'hA0;
Memory[2721] = 8'h02;
Memory[2720] = 8'h93;
Memory[2727] = 8'h02;
Memory[2726] = 8'h52;
Memory[2725] = 8'h62;
Memory[2724] = 8'h33;
Memory[2731] = 8'h00;
Memory[2730] = 8'h82;
Memory[2729] = 8'h12;
Memory[2728] = 8'h13;
Memory[2735] = 8'h00;
Memory[2734] = 8'hA0;
Memory[2733] = 8'h02;
Memory[2732] = 8'h93;
Memory[2739] = 8'h03;
Memory[2738] = 8'hB2;
Memory[2737] = 8'h82;
Memory[2736] = 8'hB3;
Memory[2743] = 8'h02;
Memory[2742] = 8'h53;
Memory[2741] = 8'hC3;
Memory[2740] = 8'h33;
Memory[2747] = 8'h00;
Memory[2746] = 8'hA0;
Memory[2745] = 8'h02;
Memory[2744] = 8'h93;
Memory[2751] = 8'h02;
Memory[2750] = 8'h53;
Memory[2749] = 8'h63;
Memory[2748] = 8'h33;
Memory[2755] = 8'h00;
Memory[2754] = 8'h62;
Memory[2753] = 8'h02;
Memory[2752] = 8'h33;
Memory[2759] = 8'h00;
Memory[2758] = 8'h41;
Memory[2757] = 8'h81;
Memory[2756] = 8'hB3;
Memory[2763] = 8'h00;
Memory[2762] = 8'h3B;
Memory[2761] = 8'h20;
Memory[2760] = 8'h23;
Memory[2767] = 8'h10;
Memory[2766] = 8'hCB;
Memory[2765] = 8'h21;
Memory[2764] = 8'h83;
Memory[2771] = 8'h3E;
Memory[2770] = 8'h80;
Memory[2769] = 8'h02;
Memory[2768] = 8'h93;
Memory[2775] = 8'h02;
Memory[2774] = 8'h53;
Memory[2773] = 8'hC2;
Memory[2772] = 8'h33;
Memory[2779] = 8'h00;
Memory[2778] = 8'hA0;
Memory[2777] = 8'h02;
Memory[2776] = 8'h93;
Memory[2783] = 8'h02;
Memory[2782] = 8'h52;
Memory[2781] = 8'h62;
Memory[2780] = 8'h33;
Memory[2787] = 8'h00;
Memory[2786] = 8'h82;
Memory[2785] = 8'h12;
Memory[2784] = 8'h13;
Memory[2791] = 8'h06;
Memory[2790] = 8'h40;
Memory[2789] = 8'h02;
Memory[2788] = 8'h93;
Memory[2795] = 8'h02;
Memory[2794] = 8'h53;
Memory[2793] = 8'hC3;
Memory[2792] = 8'h33;
Memory[2799] = 8'h00;
Memory[2798] = 8'hA0;
Memory[2797] = 8'h02;
Memory[2796] = 8'h93;
Memory[2803] = 8'h02;
Memory[2802] = 8'h53;
Memory[2801] = 8'h63;
Memory[2800] = 8'h33;
Memory[2807] = 8'h00;
Memory[2806] = 8'h62;
Memory[2805] = 8'h02;
Memory[2804] = 8'h33;
Memory[2811] = 8'h00;
Memory[2810] = 8'h82;
Memory[2809] = 8'h12;
Memory[2808] = 8'h13;
Memory[2815] = 8'h02;
Memory[2814] = 8'h53;
Memory[2813] = 8'hC3;
Memory[2812] = 8'h33;
Memory[2819] = 8'h02;
Memory[2818] = 8'h53;
Memory[2817] = 8'h63;
Memory[2816] = 8'h33;
Memory[2823] = 8'h00;
Memory[2822] = 8'h62;
Memory[2821] = 8'h02;
Memory[2820] = 8'h33;
Memory[2827] = 8'h00;
Memory[2826] = 8'h82;
Memory[2825] = 8'h12;
Memory[2824] = 8'h13;
Memory[2831] = 8'h02;
Memory[2830] = 8'h53;
Memory[2829] = 8'hE3;
Memory[2828] = 8'h33;
Memory[2835] = 8'h00;
Memory[2834] = 8'h62;
Memory[2833] = 8'h02;
Memory[2832] = 8'h33;
Memory[2839] = 8'h00;
Memory[2838] = 8'h41;
Memory[2837] = 8'h81;
Memory[2836] = 8'hB3;
Memory[2843] = 8'h00;
Memory[2842] = 8'h3B;
Memory[2841] = 8'h22;
Memory[2840] = 8'h23;
Memory[2847] = 8'h01;
Memory[2846] = 8'hDE;
Memory[2845] = 8'h14;
Memory[2844] = 8'h63;
Memory[2851] = 8'h09;
Memory[2850] = 8'hC0;
Memory[2849] = 8'h00;
Memory[2848] = 8'h6F;
Memory[2855] = 8'h01;
Memory[2854] = 8'hDE;
Memory[2853] = 8'h42;
Memory[2852] = 8'h33;
Memory[2859] = 8'h01;
Memory[2858] = 8'h82;
Memory[2857] = 8'h71;
Memory[2856] = 8'hB3;
Memory[2863] = 8'h01;
Memory[2862] = 8'hD1;
Memory[2861] = 8'hF1;
Memory[2860] = 8'hB3;
Memory[2867] = 8'h00;
Memory[2866] = 8'h01;
Memory[2865] = 8'h84;
Memory[2864] = 8'h63;
Memory[2871] = 8'h0D;
Memory[2870] = 8'h00;
Memory[2869] = 8'h20;
Memory[2868] = 8'h6F;
Memory[2875] = 8'hFF;
Memory[2874] = 8'hF2;
Memory[2873] = 8'h71;
Memory[2872] = 8'h93;
Memory[2879] = 8'h01;
Memory[2878] = 8'hD1;
Memory[2877] = 8'hF1;
Memory[2876] = 8'hB3;
Memory[2883] = 8'h00;
Memory[2882] = 8'h01;
Memory[2881] = 8'h94;
Memory[2880] = 8'h63;
Memory[2887] = 8'h2C;
Memory[2886] = 8'h40;
Memory[2885] = 8'h00;
Memory[2884] = 8'h6F;
Memory[2891] = 8'h10;
Memory[2890] = 8'h01;
Memory[2889] = 8'hF2;
Memory[2888] = 8'h13;
Memory[2895] = 8'h00;
Memory[2894] = 8'h02;
Memory[2893] = 8'h18;
Memory[2892] = 8'h63;
Memory[2899] = 8'h00;
Memory[2898] = 8'h11;
Memory[2897] = 8'hF2;
Memory[2896] = 8'h13;
Memory[2903] = 8'h00;
Memory[2902] = 8'h02;
Memory[2901] = 8'h1A;
Memory[2900] = 8'h63;
Memory[2907] = 8'h2C;
Memory[2906] = 8'h40;
Memory[2905] = 8'h00;
Memory[2904] = 8'h6F;
Memory[2911] = 8'h00;
Memory[2910] = 8'hC0;
Memory[2909] = 8'h01;
Memory[2908] = 8'h13;
Memory[2915] = 8'h00;
Memory[2914] = 8'h0E;
Memory[2913] = 8'h8E;
Memory[2912] = 8'h13;
Memory[2919] = 8'h18;
Memory[2918] = 8'h90;
Memory[2917] = 8'h00;
Memory[2916] = 8'h6F;
Memory[2923] = 8'h00;
Memory[2922] = 8'h90;
Memory[2921] = 8'h01;
Memory[2920] = 8'h13;
Memory[2927] = 8'h00;
Memory[2926] = 8'h0E;
Memory[2925] = 8'h8E;
Memory[2924] = 8'h13;
Memory[2931] = 8'h71;
Memory[2930] = 8'h80;
Memory[2929] = 8'h00;
Memory[2928] = 8'h6F;
Memory[2935] = 8'h01;
Memory[2934] = 8'h30;
Memory[2933] = 8'h01;
Memory[2932] = 8'h13;
Memory[2939] = 8'h13;
Memory[2938] = 8'h8B;
Memory[2937] = 8'h21;
Memory[2936] = 8'h83;
Memory[2943] = 8'h13;
Memory[2942] = 8'hCB;
Memory[2941] = 8'h22;
Memory[2940] = 8'h03;
Memory[2947] = 8'h00;
Memory[2946] = 8'hF0;
Memory[2945] = 8'h02;
Memory[2944] = 8'h93;
Memory[2951] = 8'h00;
Memory[2950] = 8'h3B;
Memory[2949] = 8'h20;
Memory[2948] = 8'h23;
Memory[2955] = 8'h00;
Memory[2954] = 8'h4B;
Memory[2953] = 8'h22;
Memory[2952] = 8'h23;
Memory[2959] = 8'h00;
Memory[2958] = 8'h5B;
Memory[2957] = 8'h24;
Memory[2956] = 8'h23;
Memory[2963] = 8'h01;
Memory[2962] = 8'hDE;
Memory[2961] = 8'h14;
Memory[2960] = 8'h63;
Memory[2967] = 8'h09;
Memory[2966] = 8'hC0;
Memory[2965] = 8'h00;
Memory[2964] = 8'h6F;
Memory[2971] = 8'h01;
Memory[2970] = 8'hDE;
Memory[2969] = 8'h42;
Memory[2968] = 8'h33;
Memory[2975] = 8'h01;
Memory[2974] = 8'h82;
Memory[2973] = 8'h71;
Memory[2972] = 8'hB3;
Memory[2979] = 8'h01;
Memory[2978] = 8'hD1;
Memory[2977] = 8'hF1;
Memory[2976] = 8'hB3;
Memory[2983] = 8'h00;
Memory[2982] = 8'h01;
Memory[2981] = 8'h84;
Memory[2980] = 8'h63;
Memory[2987] = 8'h0D;
Memory[2986] = 8'h00;
Memory[2985] = 8'h20;
Memory[2984] = 8'h6F;
Memory[2991] = 8'hFF;
Memory[2990] = 8'hF2;
Memory[2989] = 8'h71;
Memory[2988] = 8'h93;
Memory[2995] = 8'h01;
Memory[2994] = 8'hD1;
Memory[2993] = 8'hF1;
Memory[2992] = 8'hB3;
Memory[2999] = 8'h00;
Memory[2998] = 8'h01;
Memory[2997] = 8'h94;
Memory[2996] = 8'h63;
Memory[3003] = 8'h2C;
Memory[3002] = 8'h40;
Memory[3001] = 8'h00;
Memory[3000] = 8'h6F;
Memory[3007] = 8'h10;
Memory[3006] = 8'h01;
Memory[3005] = 8'hF2;
Memory[3004] = 8'h13;
Memory[3011] = 8'h00;
Memory[3010] = 8'h02;
Memory[3009] = 8'h1C;
Memory[3008] = 8'h63;
Memory[3015] = 8'h04;
Memory[3014] = 8'h01;
Memory[3013] = 8'hF2;
Memory[3012] = 8'h13;
Memory[3019] = 8'h00;
Memory[3018] = 8'h02;
Memory[3017] = 8'h1E;
Memory[3016] = 8'h63;
Memory[3023] = 8'h00;
Memory[3022] = 8'h41;
Memory[3021] = 8'hF2;
Memory[3020] = 8'h13;
Memory[3027] = 8'h02;
Memory[3026] = 8'h02;
Memory[3025] = 8'h10;
Memory[3024] = 8'h63;
Memory[3031] = 8'h2C;
Memory[3030] = 8'h40;
Memory[3029] = 8'h00;
Memory[3028] = 8'h6F;
Memory[3035] = 8'h00;
Memory[3034] = 8'h90;
Memory[3033] = 8'h01;
Memory[3032] = 8'h13;
Memory[3039] = 8'h00;
Memory[3038] = 8'h0E;
Memory[3037] = 8'h8E;
Memory[3036] = 8'h13;
Memory[3043] = 8'h71;
Memory[3042] = 8'h80;
Memory[3041] = 8'h00;
Memory[3040] = 8'h6F;
Memory[3047] = 8'h01;
Memory[3046] = 8'h40;
Memory[3045] = 8'h01;
Memory[3044] = 8'h13;
Memory[3051] = 8'h00;
Memory[3050] = 8'h0E;
Memory[3049] = 8'h8E;
Memory[3048] = 8'h13;
Memory[3055] = 8'h7D;
Memory[3054] = 8'h50;
Memory[3053] = 8'h00;
Memory[3052] = 8'h6F;
Memory[3059] = 8'h01;
Memory[3058] = 8'hC0;
Memory[3057] = 8'h01;
Memory[3056] = 8'h13;
Memory[3063] = 8'h00;
Memory[3062] = 8'h0E;
Memory[3061] = 8'h8E;
Memory[3060] = 8'h13;
Memory[3067] = 8'h3F;
Memory[3066] = 8'hD0;
Memory[3065] = 8'h00;
Memory[3064] = 8'h6F;
Memory[3071] = 8'h01;
Memory[3070] = 8'h40;
Memory[3069] = 8'h01;
Memory[3068] = 8'h13;
Memory[3075] = 8'h14;
Memory[3074] = 8'h0B;
Memory[3073] = 8'h21;
Memory[3072] = 8'h83;
Memory[3079] = 8'h14;
Memory[3078] = 8'h4B;
Memory[3077] = 8'h22;
Memory[3076] = 8'h03;
Memory[3083] = 8'h00;
Memory[3082] = 8'h3B;
Memory[3081] = 8'h20;
Memory[3080] = 8'h23;
Memory[3087] = 8'h00;
Memory[3086] = 8'h4B;
Memory[3085] = 8'h22;
Memory[3084] = 8'h23;
Memory[3091] = 8'h01;
Memory[3090] = 8'hDE;
Memory[3089] = 8'h14;
Memory[3088] = 8'h63;
Memory[3095] = 8'h09;
Memory[3094] = 8'hC0;
Memory[3093] = 8'h00;
Memory[3092] = 8'h6F;
Memory[3099] = 8'h01;
Memory[3098] = 8'hDE;
Memory[3097] = 8'h42;
Memory[3096] = 8'h33;
Memory[3103] = 8'h01;
Memory[3102] = 8'h82;
Memory[3101] = 8'h71;
Memory[3100] = 8'hB3;
Memory[3107] = 8'h01;
Memory[3106] = 8'hD1;
Memory[3105] = 8'hF1;
Memory[3104] = 8'hB3;
Memory[3111] = 8'h00;
Memory[3110] = 8'h01;
Memory[3109] = 8'h84;
Memory[3108] = 8'h63;
Memory[3115] = 8'h0D;
Memory[3114] = 8'h00;
Memory[3113] = 8'h20;
Memory[3112] = 8'h6F;
Memory[3119] = 8'hFF;
Memory[3118] = 8'hF2;
Memory[3117] = 8'h71;
Memory[3116] = 8'h93;
Memory[3123] = 8'h01;
Memory[3122] = 8'hD1;
Memory[3121] = 8'hF1;
Memory[3120] = 8'hB3;
Memory[3127] = 8'h00;
Memory[3126] = 8'h01;
Memory[3125] = 8'h94;
Memory[3124] = 8'h63;
Memory[3131] = 8'h2C;
Memory[3130] = 8'h40;
Memory[3129] = 8'h00;
Memory[3128] = 8'h6F;
Memory[3135] = 8'h04;
Memory[3134] = 8'h01;
Memory[3133] = 8'hF2;
Memory[3132] = 8'h13;
Memory[3139] = 8'h00;
Memory[3138] = 8'h02;
Memory[3137] = 8'h18;
Memory[3136] = 8'h63;
Memory[3143] = 8'h00;
Memory[3142] = 8'h11;
Memory[3141] = 8'hF2;
Memory[3140] = 8'h13;
Memory[3147] = 8'h00;
Memory[3146] = 8'h02;
Memory[3145] = 8'h1A;
Memory[3144] = 8'h63;
Memory[3151] = 8'h2C;
Memory[3150] = 8'h40;
Memory[3149] = 8'h00;
Memory[3148] = 8'h6F;
Memory[3155] = 8'h01;
Memory[3154] = 8'h50;
Memory[3153] = 8'h01;
Memory[3152] = 8'h13;
Memory[3159] = 8'h00;
Memory[3158] = 8'h0E;
Memory[3157] = 8'h8E;
Memory[3156] = 8'h13;
Memory[3163] = 8'h46;
Memory[3162] = 8'h90;
Memory[3161] = 8'h00;
Memory[3160] = 8'h6F;
Memory[3167] = 8'h01;
Memory[3166] = 8'h30;
Memory[3165] = 8'h01;
Memory[3164] = 8'h13;
Memory[3171] = 8'h00;
Memory[3170] = 8'h0E;
Memory[3169] = 8'h8E;
Memory[3168] = 8'h13;
Memory[3175] = 8'h37;
Memory[3174] = 8'h50;
Memory[3173] = 8'h00;
Memory[3172] = 8'h6F;
Memory[3179] = 8'h01;
Memory[3178] = 8'h50;
Memory[3177] = 8'h01;
Memory[3176] = 8'h13;
Memory[3183] = 8'h14;
Memory[3182] = 8'h8B;
Memory[3181] = 8'h21;
Memory[3180] = 8'h83;
Memory[3187] = 8'h14;
Memory[3186] = 8'hCB;
Memory[3185] = 8'h22;
Memory[3184] = 8'h03;
Memory[3191] = 8'h00;
Memory[3190] = 8'h3B;
Memory[3189] = 8'h20;
Memory[3188] = 8'h23;
Memory[3195] = 8'h00;
Memory[3194] = 8'h4B;
Memory[3193] = 8'h22;
Memory[3192] = 8'h23;
Memory[3199] = 8'h01;
Memory[3198] = 8'hDE;
Memory[3197] = 8'h14;
Memory[3196] = 8'h63;
Memory[3203] = 8'h09;
Memory[3202] = 8'hC0;
Memory[3201] = 8'h00;
Memory[3200] = 8'h6F;
Memory[3207] = 8'h01;
Memory[3206] = 8'hDE;
Memory[3205] = 8'h42;
Memory[3204] = 8'h33;
Memory[3211] = 8'h01;
Memory[3210] = 8'h82;
Memory[3209] = 8'h71;
Memory[3208] = 8'hB3;
Memory[3215] = 8'h01;
Memory[3214] = 8'hD1;
Memory[3213] = 8'hF1;
Memory[3212] = 8'hB3;
Memory[3219] = 8'h00;
Memory[3218] = 8'h01;
Memory[3217] = 8'h84;
Memory[3216] = 8'h63;
Memory[3223] = 8'h0D;
Memory[3222] = 8'h00;
Memory[3221] = 8'h20;
Memory[3220] = 8'h6F;
Memory[3227] = 8'hFF;
Memory[3226] = 8'hF2;
Memory[3225] = 8'h71;
Memory[3224] = 8'h93;
Memory[3231] = 8'h01;
Memory[3230] = 8'hD1;
Memory[3229] = 8'hF1;
Memory[3228] = 8'hB3;
Memory[3235] = 8'h00;
Memory[3234] = 8'h01;
Memory[3233] = 8'h94;
Memory[3232] = 8'h63;
Memory[3239] = 8'h2C;
Memory[3238] = 8'h40;
Memory[3237] = 8'h00;
Memory[3236] = 8'h6F;
Memory[3243] = 8'h10;
Memory[3242] = 8'h01;
Memory[3241] = 8'hF2;
Memory[3240] = 8'h13;
Memory[3247] = 8'h00;
Memory[3246] = 8'h02;
Memory[3245] = 8'h1C;
Memory[3244] = 8'h63;
Memory[3251] = 8'h04;
Memory[3250] = 8'h01;
Memory[3249] = 8'hF2;
Memory[3248] = 8'h13;
Memory[3255] = 8'h00;
Memory[3254] = 8'h02;
Memory[3253] = 8'h1E;
Memory[3252] = 8'h63;
Memory[3259] = 8'h00;
Memory[3258] = 8'h11;
Memory[3257] = 8'hF2;
Memory[3256] = 8'h13;
Memory[3263] = 8'h02;
Memory[3262] = 8'h02;
Memory[3261] = 8'h10;
Memory[3260] = 8'h63;
Memory[3267] = 8'h2C;
Memory[3266] = 8'h40;
Memory[3265] = 8'h00;
Memory[3264] = 8'h6F;
Memory[3271] = 8'h01;
Memory[3270] = 8'h40;
Memory[3269] = 8'h01;
Memory[3268] = 8'h13;
Memory[3275] = 8'h00;
Memory[3274] = 8'h0E;
Memory[3273] = 8'h8E;
Memory[3272] = 8'h13;
Memory[3279] = 8'h3F;
Memory[3278] = 8'hD0;
Memory[3277] = 8'h00;
Memory[3276] = 8'h6F;
Memory[3283] = 8'h01;
Memory[3282] = 8'h60;
Memory[3281] = 8'h01;
Memory[3280] = 8'h13;
Memory[3287] = 8'h00;
Memory[3286] = 8'h0E;
Memory[3285] = 8'h8E;
Memory[3284] = 8'h13;
Memory[3291] = 8'h4E;
Memory[3290] = 8'h90;
Memory[3289] = 8'h00;
Memory[3288] = 8'h6F;
Memory[3295] = 8'h01;
Memory[3294] = 8'h30;
Memory[3293] = 8'h01;
Memory[3292] = 8'h13;
Memory[3299] = 8'h00;
Memory[3298] = 8'h0E;
Memory[3297] = 8'h8E;
Memory[3296] = 8'h13;
Memory[3303] = 8'h37;
Memory[3302] = 8'h50;
Memory[3301] = 8'h00;
Memory[3300] = 8'h6F;
Memory[3307] = 8'h01;
Memory[3306] = 8'h60;
Memory[3305] = 8'h01;
Memory[3304] = 8'h13;
Memory[3311] = 8'h15;
Memory[3310] = 8'h0B;
Memory[3309] = 8'h21;
Memory[3308] = 8'h83;
Memory[3315] = 8'h15;
Memory[3314] = 8'h4B;
Memory[3313] = 8'h22;
Memory[3312] = 8'h03;
Memory[3319] = 8'h00;
Memory[3318] = 8'h3B;
Memory[3317] = 8'h20;
Memory[3316] = 8'h23;
Memory[3323] = 8'h00;
Memory[3322] = 8'h4B;
Memory[3321] = 8'h22;
Memory[3320] = 8'h23;
Memory[3327] = 8'h01;
Memory[3326] = 8'hDE;
Memory[3325] = 8'h14;
Memory[3324] = 8'h63;
Memory[3331] = 8'h09;
Memory[3330] = 8'hC0;
Memory[3329] = 8'h00;
Memory[3328] = 8'h6F;
Memory[3335] = 8'h01;
Memory[3334] = 8'hDE;
Memory[3333] = 8'h42;
Memory[3332] = 8'h33;
Memory[3339] = 8'h01;
Memory[3338] = 8'h82;
Memory[3337] = 8'h71;
Memory[3336] = 8'hB3;
Memory[3343] = 8'h01;
Memory[3342] = 8'hD1;
Memory[3341] = 8'hF1;
Memory[3340] = 8'hB3;
Memory[3347] = 8'h00;
Memory[3346] = 8'h01;
Memory[3345] = 8'h84;
Memory[3344] = 8'h63;
Memory[3351] = 8'h0D;
Memory[3350] = 8'h00;
Memory[3349] = 8'h20;
Memory[3348] = 8'h6F;
Memory[3355] = 8'hFF;
Memory[3354] = 8'hF2;
Memory[3353] = 8'h71;
Memory[3352] = 8'h93;
Memory[3359] = 8'h01;
Memory[3358] = 8'hD1;
Memory[3357] = 8'hF1;
Memory[3356] = 8'hB3;
Memory[3363] = 8'h00;
Memory[3362] = 8'h01;
Memory[3361] = 8'h94;
Memory[3360] = 8'h63;
Memory[3367] = 8'h2C;
Memory[3366] = 8'h40;
Memory[3365] = 8'h00;
Memory[3364] = 8'h6F;
Memory[3371] = 8'h10;
Memory[3370] = 8'h01;
Memory[3369] = 8'hF2;
Memory[3368] = 8'h13;
Memory[3375] = 8'h00;
Memory[3374] = 8'h02;
Memory[3373] = 8'h1C;
Memory[3372] = 8'h63;
Memory[3379] = 8'h04;
Memory[3378] = 8'h01;
Memory[3377] = 8'hF2;
Memory[3376] = 8'h13;
Memory[3383] = 8'h00;
Memory[3382] = 8'h02;
Memory[3381] = 8'h1E;
Memory[3380] = 8'h63;
Memory[3387] = 8'h00;
Memory[3386] = 8'h11;
Memory[3385] = 8'hF2;
Memory[3384] = 8'h13;
Memory[3391] = 8'h02;
Memory[3390] = 8'h02;
Memory[3389] = 8'h10;
Memory[3388] = 8'h63;
Memory[3395] = 8'h2C;
Memory[3394] = 8'h40;
Memory[3393] = 8'h00;
Memory[3392] = 8'h6F;
Memory[3399] = 8'h01;
Memory[3398] = 8'h50;
Memory[3397] = 8'h01;
Memory[3396] = 8'h13;
Memory[3403] = 8'h00;
Memory[3402] = 8'h0E;
Memory[3401] = 8'h8E;
Memory[3400] = 8'h13;
Memory[3407] = 8'h46;
Memory[3406] = 8'h90;
Memory[3405] = 8'h00;
Memory[3404] = 8'h6F;
Memory[3411] = 8'h01;
Memory[3410] = 8'h70;
Memory[3409] = 8'h01;
Memory[3408] = 8'h13;
Memory[3415] = 8'h00;
Memory[3414] = 8'h0E;
Memory[3413] = 8'h8E;
Memory[3412] = 8'h13;
Memory[3419] = 8'h56;
Memory[3418] = 8'h90;
Memory[3417] = 8'h00;
Memory[3416] = 8'h6F;
Memory[3423] = 8'h01;
Memory[3422] = 8'h30;
Memory[3421] = 8'h01;
Memory[3420] = 8'h13;
Memory[3427] = 8'h00;
Memory[3426] = 8'h0E;
Memory[3425] = 8'h8E;
Memory[3424] = 8'h13;
Memory[3431] = 8'h37;
Memory[3430] = 8'h50;
Memory[3429] = 8'h00;
Memory[3428] = 8'h6F;
Memory[3435] = 8'h01;
Memory[3434] = 8'h70;
Memory[3433] = 8'h01;
Memory[3432] = 8'h13;
Memory[3439] = 8'h15;
Memory[3438] = 8'h8B;
Memory[3437] = 8'h21;
Memory[3436] = 8'h83;
Memory[3443] = 8'h15;
Memory[3442] = 8'hCB;
Memory[3441] = 8'h22;
Memory[3440] = 8'h03;
Memory[3447] = 8'h00;
Memory[3446] = 8'h3B;
Memory[3445] = 8'h20;
Memory[3444] = 8'h23;
Memory[3451] = 8'h00;
Memory[3450] = 8'h4B;
Memory[3449] = 8'h22;
Memory[3448] = 8'h23;
Memory[3455] = 8'h01;
Memory[3454] = 8'hDE;
Memory[3453] = 8'h14;
Memory[3452] = 8'h63;
Memory[3459] = 8'h09;
Memory[3458] = 8'hC0;
Memory[3457] = 8'h00;
Memory[3456] = 8'h6F;
Memory[3463] = 8'h01;
Memory[3462] = 8'hDE;
Memory[3461] = 8'h42;
Memory[3460] = 8'h33;
Memory[3467] = 8'h01;
Memory[3466] = 8'h82;
Memory[3465] = 8'h71;
Memory[3464] = 8'hB3;
Memory[3471] = 8'h01;
Memory[3470] = 8'hD1;
Memory[3469] = 8'hF1;
Memory[3468] = 8'hB3;
Memory[3475] = 8'h00;
Memory[3474] = 8'h01;
Memory[3473] = 8'h84;
Memory[3472] = 8'h63;
Memory[3479] = 8'h0D;
Memory[3478] = 8'h00;
Memory[3477] = 8'h20;
Memory[3476] = 8'h6F;
Memory[3483] = 8'hFF;
Memory[3482] = 8'hF2;
Memory[3481] = 8'h71;
Memory[3480] = 8'h93;
Memory[3487] = 8'h01;
Memory[3486] = 8'hD1;
Memory[3485] = 8'hF1;
Memory[3484] = 8'hB3;
Memory[3491] = 8'h00;
Memory[3490] = 8'h01;
Memory[3489] = 8'h94;
Memory[3488] = 8'h63;
Memory[3495] = 8'h2C;
Memory[3494] = 8'h40;
Memory[3493] = 8'h00;
Memory[3492] = 8'h6F;
Memory[3499] = 8'h10;
Memory[3498] = 8'h01;
Memory[3497] = 8'hF2;
Memory[3496] = 8'h13;
Memory[3503] = 8'h00;
Memory[3502] = 8'h02;
Memory[3501] = 8'h1C;
Memory[3500] = 8'h63;
Memory[3507] = 8'h04;
Memory[3506] = 8'h01;
Memory[3505] = 8'hF2;
Memory[3504] = 8'h13;
Memory[3511] = 8'h00;
Memory[3510] = 8'h02;
Memory[3509] = 8'h1E;
Memory[3508] = 8'h63;
Memory[3515] = 8'h00;
Memory[3514] = 8'h11;
Memory[3513] = 8'hF2;
Memory[3512] = 8'h13;
Memory[3519] = 8'h02;
Memory[3518] = 8'h02;
Memory[3517] = 8'h10;
Memory[3516] = 8'h63;
Memory[3523] = 8'h2C;
Memory[3522] = 8'h40;
Memory[3521] = 8'h00;
Memory[3520] = 8'h6F;
Memory[3527] = 8'h01;
Memory[3526] = 8'h60;
Memory[3525] = 8'h01;
Memory[3524] = 8'h13;
Memory[3531] = 8'h00;
Memory[3530] = 8'h0E;
Memory[3529] = 8'h8E;
Memory[3528] = 8'h13;
Memory[3535] = 8'h4E;
Memory[3534] = 8'h90;
Memory[3533] = 8'h00;
Memory[3532] = 8'h6F;
Memory[3539] = 8'h01;
Memory[3538] = 8'h80;
Memory[3537] = 8'h01;
Memory[3536] = 8'h13;
Memory[3543] = 8'h00;
Memory[3542] = 8'h0E;
Memory[3541] = 8'h8E;
Memory[3540] = 8'h13;
Memory[3547] = 8'h5E;
Memory[3546] = 8'h90;
Memory[3545] = 8'h00;
Memory[3544] = 8'h6F;
Memory[3551] = 8'h01;
Memory[3550] = 8'h30;
Memory[3549] = 8'h01;
Memory[3548] = 8'h13;
Memory[3555] = 8'h00;
Memory[3554] = 8'h0E;
Memory[3553] = 8'h8E;
Memory[3552] = 8'h13;
Memory[3559] = 8'h37;
Memory[3558] = 8'h50;
Memory[3557] = 8'h00;
Memory[3556] = 8'h6F;
Memory[3563] = 8'h01;
Memory[3562] = 8'h80;
Memory[3561] = 8'h01;
Memory[3560] = 8'h13;
Memory[3567] = 8'h16;
Memory[3566] = 8'h0B;
Memory[3565] = 8'h21;
Memory[3564] = 8'h83;
Memory[3571] = 8'h16;
Memory[3570] = 8'h4B;
Memory[3569] = 8'h22;
Memory[3568] = 8'h03;
Memory[3575] = 8'h00;
Memory[3574] = 8'h3B;
Memory[3573] = 8'h20;
Memory[3572] = 8'h23;
Memory[3579] = 8'h00;
Memory[3578] = 8'h4B;
Memory[3577] = 8'h22;
Memory[3576] = 8'h23;
Memory[3583] = 8'h01;
Memory[3582] = 8'hDE;
Memory[3581] = 8'h14;
Memory[3580] = 8'h63;
Memory[3587] = 8'h09;
Memory[3586] = 8'hC0;
Memory[3585] = 8'h00;
Memory[3584] = 8'h6F;
Memory[3591] = 8'h01;
Memory[3590] = 8'hDE;
Memory[3589] = 8'h42;
Memory[3588] = 8'h33;
Memory[3595] = 8'h01;
Memory[3594] = 8'h82;
Memory[3593] = 8'h71;
Memory[3592] = 8'hB3;
Memory[3599] = 8'h01;
Memory[3598] = 8'hD1;
Memory[3597] = 8'hF1;
Memory[3596] = 8'hB3;
Memory[3603] = 8'h00;
Memory[3602] = 8'h01;
Memory[3601] = 8'h84;
Memory[3600] = 8'h63;
Memory[3607] = 8'h0D;
Memory[3606] = 8'h00;
Memory[3605] = 8'h20;
Memory[3604] = 8'h6F;
Memory[3611] = 8'hFF;
Memory[3610] = 8'hF2;
Memory[3609] = 8'h71;
Memory[3608] = 8'h93;
Memory[3615] = 8'h01;
Memory[3614] = 8'hD1;
Memory[3613] = 8'hF1;
Memory[3612] = 8'hB3;
Memory[3619] = 8'h00;
Memory[3618] = 8'h01;
Memory[3617] = 8'h94;
Memory[3616] = 8'h63;
Memory[3623] = 8'h2C;
Memory[3622] = 8'h40;
Memory[3621] = 8'h00;
Memory[3620] = 8'h6F;
Memory[3627] = 8'h10;
Memory[3626] = 8'h01;
Memory[3625] = 8'hF2;
Memory[3624] = 8'h13;
Memory[3631] = 8'h00;
Memory[3630] = 8'h02;
Memory[3629] = 8'h1C;
Memory[3628] = 8'h63;
Memory[3635] = 8'h04;
Memory[3634] = 8'h01;
Memory[3633] = 8'hF2;
Memory[3632] = 8'h13;
Memory[3639] = 8'h00;
Memory[3638] = 8'h02;
Memory[3637] = 8'h1E;
Memory[3636] = 8'h63;
Memory[3643] = 8'h00;
Memory[3642] = 8'h11;
Memory[3641] = 8'hF2;
Memory[3640] = 8'h13;
Memory[3647] = 8'h02;
Memory[3646] = 8'h02;
Memory[3645] = 8'h10;
Memory[3644] = 8'h63;
Memory[3651] = 8'h2C;
Memory[3650] = 8'h40;
Memory[3649] = 8'h00;
Memory[3648] = 8'h6F;
Memory[3655] = 8'h01;
Memory[3654] = 8'h70;
Memory[3653] = 8'h01;
Memory[3652] = 8'h13;
Memory[3659] = 8'h00;
Memory[3658] = 8'h0E;
Memory[3657] = 8'h8E;
Memory[3656] = 8'h13;
Memory[3663] = 8'h56;
Memory[3662] = 8'h90;
Memory[3661] = 8'h00;
Memory[3660] = 8'h6F;
Memory[3667] = 8'h01;
Memory[3666] = 8'h90;
Memory[3665] = 8'h01;
Memory[3664] = 8'h13;
Memory[3671] = 8'h00;
Memory[3670] = 8'h0E;
Memory[3669] = 8'h8E;
Memory[3668] = 8'h13;
Memory[3675] = 8'h66;
Memory[3674] = 8'h90;
Memory[3673] = 8'h00;
Memory[3672] = 8'h6F;
Memory[3679] = 8'h01;
Memory[3678] = 8'h30;
Memory[3677] = 8'h01;
Memory[3676] = 8'h13;
Memory[3683] = 8'h00;
Memory[3682] = 8'h0E;
Memory[3681] = 8'h8E;
Memory[3680] = 8'h13;
Memory[3687] = 8'h37;
Memory[3686] = 8'h50;
Memory[3685] = 8'h00;
Memory[3684] = 8'h6F;
Memory[3691] = 8'h01;
Memory[3690] = 8'h90;
Memory[3689] = 8'h01;
Memory[3688] = 8'h13;
Memory[3695] = 8'h16;
Memory[3694] = 8'h8B;
Memory[3693] = 8'h21;
Memory[3692] = 8'h83;
Memory[3699] = 8'h16;
Memory[3698] = 8'hCB;
Memory[3697] = 8'h22;
Memory[3696] = 8'h03;
Memory[3703] = 8'h00;
Memory[3702] = 8'h3B;
Memory[3701] = 8'h20;
Memory[3700] = 8'h23;
Memory[3707] = 8'h00;
Memory[3706] = 8'h4B;
Memory[3705] = 8'h22;
Memory[3704] = 8'h23;
Memory[3711] = 8'h01;
Memory[3710] = 8'hDE;
Memory[3709] = 8'h14;
Memory[3708] = 8'h63;
Memory[3715] = 8'h09;
Memory[3714] = 8'hC0;
Memory[3713] = 8'h00;
Memory[3712] = 8'h6F;
Memory[3719] = 8'h01;
Memory[3718] = 8'hDE;
Memory[3717] = 8'h42;
Memory[3716] = 8'h33;
Memory[3723] = 8'h01;
Memory[3722] = 8'h82;
Memory[3721] = 8'h71;
Memory[3720] = 8'hB3;
Memory[3727] = 8'h01;
Memory[3726] = 8'hD1;
Memory[3725] = 8'hF1;
Memory[3724] = 8'hB3;
Memory[3731] = 8'h00;
Memory[3730] = 8'h01;
Memory[3729] = 8'h84;
Memory[3728] = 8'h63;
Memory[3735] = 8'h0D;
Memory[3734] = 8'h00;
Memory[3733] = 8'h20;
Memory[3732] = 8'h6F;
Memory[3739] = 8'hFF;
Memory[3738] = 8'hF2;
Memory[3737] = 8'h71;
Memory[3736] = 8'h93;
Memory[3743] = 8'h01;
Memory[3742] = 8'hD1;
Memory[3741] = 8'hF1;
Memory[3740] = 8'hB3;
Memory[3747] = 8'h00;
Memory[3746] = 8'h01;
Memory[3745] = 8'h94;
Memory[3744] = 8'h63;
Memory[3751] = 8'h2C;
Memory[3750] = 8'h40;
Memory[3749] = 8'h00;
Memory[3748] = 8'h6F;
Memory[3755] = 8'h10;
Memory[3754] = 8'h01;
Memory[3753] = 8'hF2;
Memory[3752] = 8'h13;
Memory[3759] = 8'h00;
Memory[3758] = 8'h02;
Memory[3757] = 8'h1C;
Memory[3756] = 8'h63;
Memory[3763] = 8'h04;
Memory[3762] = 8'h01;
Memory[3761] = 8'hF2;
Memory[3760] = 8'h13;
Memory[3767] = 8'h00;
Memory[3766] = 8'h02;
Memory[3765] = 8'h1E;
Memory[3764] = 8'h63;
Memory[3771] = 8'h00;
Memory[3770] = 8'h11;
Memory[3769] = 8'hF2;
Memory[3768] = 8'h13;
Memory[3775] = 8'h02;
Memory[3774] = 8'h02;
Memory[3773] = 8'h10;
Memory[3772] = 8'h63;
Memory[3779] = 8'h2C;
Memory[3778] = 8'h40;
Memory[3777] = 8'h00;
Memory[3776] = 8'h6F;
Memory[3783] = 8'h01;
Memory[3782] = 8'h80;
Memory[3781] = 8'h01;
Memory[3780] = 8'h13;
Memory[3787] = 8'h00;
Memory[3786] = 8'h0E;
Memory[3785] = 8'h8E;
Memory[3784] = 8'h13;
Memory[3791] = 8'h5E;
Memory[3790] = 8'h90;
Memory[3789] = 8'h00;
Memory[3788] = 8'h6F;
Memory[3795] = 8'h01;
Memory[3794] = 8'hA0;
Memory[3793] = 8'h01;
Memory[3792] = 8'h13;
Memory[3799] = 8'h00;
Memory[3798] = 8'h0E;
Memory[3797] = 8'h8E;
Memory[3796] = 8'h13;
Memory[3803] = 8'h6E;
Memory[3802] = 8'h90;
Memory[3801] = 8'h00;
Memory[3800] = 8'h6F;
Memory[3807] = 8'h01;
Memory[3806] = 8'h30;
Memory[3805] = 8'h01;
Memory[3804] = 8'h13;
Memory[3811] = 8'h00;
Memory[3810] = 8'h0E;
Memory[3809] = 8'h8E;
Memory[3808] = 8'h13;
Memory[3815] = 8'h37;
Memory[3814] = 8'h50;
Memory[3813] = 8'h00;
Memory[3812] = 8'h6F;
Memory[3819] = 8'h01;
Memory[3818] = 8'hA0;
Memory[3817] = 8'h01;
Memory[3816] = 8'h13;
Memory[3823] = 8'h17;
Memory[3822] = 8'h0B;
Memory[3821] = 8'h21;
Memory[3820] = 8'h83;
Memory[3827] = 8'h17;
Memory[3826] = 8'h4B;
Memory[3825] = 8'h22;
Memory[3824] = 8'h03;
Memory[3831] = 8'h00;
Memory[3830] = 8'h3B;
Memory[3829] = 8'h20;
Memory[3828] = 8'h23;
Memory[3835] = 8'h00;
Memory[3834] = 8'h4B;
Memory[3833] = 8'h22;
Memory[3832] = 8'h23;
Memory[3839] = 8'h01;
Memory[3838] = 8'hDE;
Memory[3837] = 8'h14;
Memory[3836] = 8'h63;
Memory[3843] = 8'h09;
Memory[3842] = 8'hC0;
Memory[3841] = 8'h00;
Memory[3840] = 8'h6F;
Memory[3847] = 8'h01;
Memory[3846] = 8'hDE;
Memory[3845] = 8'h42;
Memory[3844] = 8'h33;
Memory[3851] = 8'h01;
Memory[3850] = 8'h82;
Memory[3849] = 8'h71;
Memory[3848] = 8'hB3;
Memory[3855] = 8'h01;
Memory[3854] = 8'hD1;
Memory[3853] = 8'hF1;
Memory[3852] = 8'hB3;
Memory[3859] = 8'h00;
Memory[3858] = 8'h01;
Memory[3857] = 8'h84;
Memory[3856] = 8'h63;
Memory[3863] = 8'h0D;
Memory[3862] = 8'h00;
Memory[3861] = 8'h20;
Memory[3860] = 8'h6F;
Memory[3867] = 8'hFF;
Memory[3866] = 8'hF2;
Memory[3865] = 8'h71;
Memory[3864] = 8'h93;
Memory[3871] = 8'h01;
Memory[3870] = 8'hD1;
Memory[3869] = 8'hF1;
Memory[3868] = 8'hB3;
Memory[3875] = 8'h00;
Memory[3874] = 8'h01;
Memory[3873] = 8'h94;
Memory[3872] = 8'h63;
Memory[3879] = 8'h2C;
Memory[3878] = 8'h40;
Memory[3877] = 8'h00;
Memory[3876] = 8'h6F;
Memory[3883] = 8'h10;
Memory[3882] = 8'h01;
Memory[3881] = 8'hF2;
Memory[3880] = 8'h13;
Memory[3887] = 8'h00;
Memory[3886] = 8'h02;
Memory[3885] = 8'h1C;
Memory[3884] = 8'h63;
Memory[3891] = 8'h04;
Memory[3890] = 8'h01;
Memory[3889] = 8'hF2;
Memory[3888] = 8'h13;
Memory[3895] = 8'h00;
Memory[3894] = 8'h02;
Memory[3893] = 8'h1E;
Memory[3892] = 8'h63;
Memory[3899] = 8'h00;
Memory[3898] = 8'h11;
Memory[3897] = 8'hF2;
Memory[3896] = 8'h13;
Memory[3903] = 8'h02;
Memory[3902] = 8'h02;
Memory[3901] = 8'h10;
Memory[3900] = 8'h63;
Memory[3907] = 8'h2C;
Memory[3906] = 8'h40;
Memory[3905] = 8'h00;
Memory[3904] = 8'h6F;
Memory[3911] = 8'h01;
Memory[3910] = 8'h90;
Memory[3909] = 8'h01;
Memory[3908] = 8'h13;
Memory[3915] = 8'h00;
Memory[3914] = 8'h0E;
Memory[3913] = 8'h8E;
Memory[3912] = 8'h13;
Memory[3919] = 8'h66;
Memory[3918] = 8'h90;
Memory[3917] = 8'h00;
Memory[3916] = 8'h6F;
Memory[3923] = 8'h01;
Memory[3922] = 8'hB0;
Memory[3921] = 8'h01;
Memory[3920] = 8'h13;
Memory[3927] = 8'h00;
Memory[3926] = 8'h0E;
Memory[3925] = 8'h8E;
Memory[3924] = 8'h13;
Memory[3931] = 8'h76;
Memory[3930] = 8'h90;
Memory[3929] = 8'h00;
Memory[3928] = 8'h6F;
Memory[3935] = 8'h01;
Memory[3934] = 8'h30;
Memory[3933] = 8'h01;
Memory[3932] = 8'h13;
Memory[3939] = 8'h00;
Memory[3938] = 8'h0E;
Memory[3937] = 8'h8E;
Memory[3936] = 8'h13;
Memory[3943] = 8'h37;
Memory[3942] = 8'h50;
Memory[3941] = 8'h00;
Memory[3940] = 8'h6F;
Memory[3947] = 8'h01;
Memory[3946] = 8'hB0;
Memory[3945] = 8'h01;
Memory[3944] = 8'h13;
Memory[3951] = 8'h17;
Memory[3950] = 8'h8B;
Memory[3949] = 8'h21;
Memory[3948] = 8'h83;
Memory[3955] = 8'h17;
Memory[3954] = 8'hCB;
Memory[3953] = 8'h22;
Memory[3952] = 8'h03;
Memory[3959] = 8'h00;
Memory[3958] = 8'h3B;
Memory[3957] = 8'h20;
Memory[3956] = 8'h23;
Memory[3963] = 8'h00;
Memory[3962] = 8'h4B;
Memory[3961] = 8'h22;
Memory[3960] = 8'h23;
Memory[3967] = 8'h01;
Memory[3966] = 8'hDE;
Memory[3965] = 8'h14;
Memory[3964] = 8'h63;
Memory[3971] = 8'h09;
Memory[3970] = 8'hC0;
Memory[3969] = 8'h00;
Memory[3968] = 8'h6F;
Memory[3975] = 8'h01;
Memory[3974] = 8'hDE;
Memory[3973] = 8'h42;
Memory[3972] = 8'h33;
Memory[3979] = 8'h01;
Memory[3978] = 8'h82;
Memory[3977] = 8'h71;
Memory[3976] = 8'hB3;
Memory[3983] = 8'h01;
Memory[3982] = 8'hD1;
Memory[3981] = 8'hF1;
Memory[3980] = 8'hB3;
Memory[3987] = 8'h00;
Memory[3986] = 8'h01;
Memory[3985] = 8'h84;
Memory[3984] = 8'h63;
Memory[3991] = 8'h0D;
Memory[3990] = 8'h00;
Memory[3989] = 8'h20;
Memory[3988] = 8'h6F;
Memory[3995] = 8'hFF;
Memory[3994] = 8'hF2;
Memory[3993] = 8'h71;
Memory[3992] = 8'h93;
Memory[3999] = 8'h01;
Memory[3998] = 8'hD1;
Memory[3997] = 8'hF1;
Memory[3996] = 8'hB3;
Memory[4003] = 8'h00;
Memory[4002] = 8'h01;
Memory[4001] = 8'h94;
Memory[4000] = 8'h63;
Memory[4007] = 8'h2C;
Memory[4006] = 8'h40;
Memory[4005] = 8'h00;
Memory[4004] = 8'h6F;
Memory[4011] = 8'h10;
Memory[4010] = 8'h01;
Memory[4009] = 8'hF2;
Memory[4008] = 8'h13;
Memory[4015] = 8'h00;
Memory[4014] = 8'h02;
Memory[4013] = 8'h18;
Memory[4012] = 8'h63;
Memory[4019] = 8'h00;
Memory[4018] = 8'h11;
Memory[4017] = 8'hF2;
Memory[4016] = 8'h13;
Memory[4023] = 8'h00;
Memory[4022] = 8'h02;
Memory[4021] = 8'h1A;
Memory[4020] = 8'h63;
Memory[4027] = 8'h2C;
Memory[4026] = 8'h40;
Memory[4025] = 8'h00;
Memory[4024] = 8'h6F;
Memory[4031] = 8'h01;
Memory[4030] = 8'hA0;
Memory[4029] = 8'h01;
Memory[4028] = 8'h13;
Memory[4035] = 8'h00;
Memory[4034] = 8'h0E;
Memory[4033] = 8'h8E;
Memory[4032] = 8'h13;
Memory[4039] = 8'h6E;
Memory[4038] = 8'h90;
Memory[4037] = 8'h00;
Memory[4036] = 8'h6F;
Memory[4043] = 8'h01;
Memory[4042] = 8'h30;
Memory[4041] = 8'h01;
Memory[4040] = 8'h13;
Memory[4047] = 8'h00;
Memory[4046] = 8'h0E;
Memory[4045] = 8'h8E;
Memory[4044] = 8'h13;
Memory[4051] = 8'h37;
Memory[4050] = 8'h50;
Memory[4049] = 8'h00;
Memory[4048] = 8'h6F;
Memory[4055] = 8'h01;
Memory[4054] = 8'hC0;
Memory[4053] = 8'h01;
Memory[4052] = 8'h13;
Memory[4059] = 8'h18;
Memory[4058] = 8'h0B;
Memory[4057] = 8'h21;
Memory[4056] = 8'h83;
Memory[4063] = 8'h18;
Memory[4062] = 8'h4B;
Memory[4061] = 8'h22;
Memory[4060] = 8'h03;
Memory[4067] = 8'h01;
Memory[4066] = 8'hB0;
Memory[4065] = 8'h02;
Memory[4064] = 8'h93;
Memory[4071] = 8'h00;
Memory[4070] = 8'h3B;
Memory[4069] = 8'h20;
Memory[4068] = 8'h23;
Memory[4075] = 8'h00;
Memory[4074] = 8'h4B;
Memory[4073] = 8'h22;
Memory[4072] = 8'h23;
Memory[4079] = 8'h00;
Memory[4078] = 8'h5B;
Memory[4077] = 8'h24;
Memory[4076] = 8'h23;
Memory[4083] = 8'h01;
Memory[4082] = 8'hDE;
Memory[4081] = 8'h14;
Memory[4080] = 8'h63;
Memory[4087] = 8'h09;
Memory[4086] = 8'hC0;
Memory[4085] = 8'h00;
Memory[4084] = 8'h6F;
Memory[4091] = 8'h01;
Memory[4090] = 8'hDE;
Memory[4089] = 8'h42;
Memory[4088] = 8'h33;
Memory[4095] = 8'h01;
Memory[4094] = 8'h82;
Memory[4093] = 8'h71;
Memory[4092] = 8'hB3;
Memory[4099] = 8'h01;
Memory[4098] = 8'hD1;
Memory[4097] = 8'hF1;
Memory[4096] = 8'hB3;
Memory[4103] = 8'h00;
Memory[4102] = 8'h01;
Memory[4101] = 8'h84;
Memory[4100] = 8'h63;
Memory[4107] = 8'h0D;
Memory[4106] = 8'h00;
Memory[4105] = 8'h20;
Memory[4104] = 8'h6F;
Memory[4111] = 8'hFF;
Memory[4110] = 8'hF2;
Memory[4109] = 8'h71;
Memory[4108] = 8'h93;
Memory[4115] = 8'h01;
Memory[4114] = 8'hD1;
Memory[4113] = 8'hF1;
Memory[4112] = 8'hB3;
Memory[4119] = 8'h00;
Memory[4118] = 8'h01;
Memory[4117] = 8'h94;
Memory[4116] = 8'h63;
Memory[4123] = 8'h2C;
Memory[4122] = 8'h40;
Memory[4121] = 8'h00;
Memory[4120] = 8'h6F;
Memory[4127] = 8'h10;
Memory[4126] = 8'h01;
Memory[4125] = 8'hF2;
Memory[4124] = 8'h13;
Memory[4131] = 8'h00;
Memory[4130] = 8'h02;
Memory[4129] = 8'h18;
Memory[4128] = 8'h63;
Memory[4135] = 8'h00;
Memory[4134] = 8'h41;
Memory[4133] = 8'hF2;
Memory[4132] = 8'h13;
Memory[4139] = 8'h00;
Memory[4138] = 8'h02;
Memory[4137] = 8'h1A;
Memory[4136] = 8'h63;
Memory[4143] = 8'h2C;
Memory[4142] = 8'h40;
Memory[4141] = 8'h00;
Memory[4140] = 8'h6F;
Memory[4147] = 8'h01;
Memory[4146] = 8'h30;
Memory[4145] = 8'h01;
Memory[4144] = 8'h13;
Memory[4151] = 8'h00;
Memory[4150] = 8'h0E;
Memory[4149] = 8'h8E;
Memory[4148] = 8'h13;
Memory[4155] = 8'h37;
Memory[4154] = 8'h50;
Memory[4153] = 8'h00;
Memory[4152] = 8'h6F;
Memory[4159] = 8'h01;
Memory[4158] = 8'hD0;
Memory[4157] = 8'h01;
Memory[4156] = 8'h13;
Memory[4163] = 8'h00;
Memory[4162] = 8'h0E;
Memory[4161] = 8'h8E;
Memory[4160] = 8'h13;
Memory[4167] = 8'h04;
Memory[4166] = 8'h80;
Memory[4165] = 8'h10;
Memory[4164] = 8'h6F;
Memory[4171] = 8'h01;
Memory[4170] = 8'hD0;
Memory[4169] = 8'h01;
Memory[4168] = 8'h13;
Memory[4175] = 8'h18;
Memory[4174] = 8'h8B;
Memory[4173] = 8'h21;
Memory[4172] = 8'h83;
Memory[4179] = 8'h18;
Memory[4178] = 8'hCB;
Memory[4177] = 8'h22;
Memory[4176] = 8'h03;
Memory[4183] = 8'h00;
Memory[4182] = 8'hB0;
Memory[4181] = 8'h02;
Memory[4180] = 8'h93;
Memory[4187] = 8'h00;
Memory[4186] = 8'h3B;
Memory[4185] = 8'h20;
Memory[4184] = 8'h23;
Memory[4191] = 8'h00;
Memory[4190] = 8'h4B;
Memory[4189] = 8'h22;
Memory[4188] = 8'h23;
Memory[4195] = 8'h00;
Memory[4194] = 8'h5B;
Memory[4193] = 8'h24;
Memory[4192] = 8'h23;
Memory[4199] = 8'h01;
Memory[4198] = 8'hDE;
Memory[4197] = 8'h14;
Memory[4196] = 8'h63;
Memory[4203] = 8'h09;
Memory[4202] = 8'hC0;
Memory[4201] = 8'h00;
Memory[4200] = 8'h6F;
Memory[4207] = 8'h01;
Memory[4206] = 8'hDE;
Memory[4205] = 8'h42;
Memory[4204] = 8'h33;
Memory[4211] = 8'h01;
Memory[4210] = 8'h82;
Memory[4209] = 8'h71;
Memory[4208] = 8'hB3;
Memory[4215] = 8'h01;
Memory[4214] = 8'hD1;
Memory[4213] = 8'hF1;
Memory[4212] = 8'hB3;
Memory[4219] = 8'h00;
Memory[4218] = 8'h01;
Memory[4217] = 8'h84;
Memory[4216] = 8'h63;
Memory[4223] = 8'h0D;
Memory[4222] = 8'h00;
Memory[4221] = 8'h20;
Memory[4220] = 8'h6F;
Memory[4227] = 8'hFF;
Memory[4226] = 8'hF2;
Memory[4225] = 8'h71;
Memory[4224] = 8'h93;
Memory[4231] = 8'h01;
Memory[4230] = 8'hD1;
Memory[4229] = 8'hF1;
Memory[4228] = 8'hB3;
Memory[4235] = 8'h00;
Memory[4234] = 8'h01;
Memory[4233] = 8'h94;
Memory[4232] = 8'h63;
Memory[4239] = 8'h2C;
Memory[4238] = 8'h40;
Memory[4237] = 8'h00;
Memory[4236] = 8'h6F;
Memory[4243] = 8'h01;
Memory[4242] = 8'h01;
Memory[4241] = 8'hF2;
Memory[4240] = 8'h13;
Memory[4247] = 8'h00;
Memory[4246] = 8'h02;
Memory[4245] = 8'h1C;
Memory[4244] = 8'h63;
Memory[4251] = 8'h00;
Memory[4250] = 8'h41;
Memory[4249] = 8'hF2;
Memory[4248] = 8'h13;
Memory[4255] = 8'h00;
Memory[4254] = 8'h02;
Memory[4253] = 8'h1E;
Memory[4252] = 8'h63;
Memory[4259] = 8'h00;
Memory[4258] = 8'h11;
Memory[4257] = 8'hF2;
Memory[4256] = 8'h13;
Memory[4263] = 8'h02;
Memory[4262] = 8'h02;
Memory[4261] = 8'h10;
Memory[4260] = 8'h63;
Memory[4267] = 8'h2C;
Memory[4266] = 8'h40;
Memory[4265] = 8'h00;
Memory[4264] = 8'h6F;
Memory[4271] = 8'h01;
Memory[4270] = 8'hF0;
Memory[4269] = 8'h01;
Memory[4268] = 8'h13;
Memory[4275] = 8'h00;
Memory[4274] = 8'h0E;
Memory[4273] = 8'h8E;
Memory[4272] = 8'h13;
Memory[4279] = 8'h32;
Memory[4278] = 8'h40;
Memory[4277] = 8'h10;
Memory[4276] = 8'h6F;
Memory[4283] = 8'h01;
Memory[4282] = 8'hE0;
Memory[4281] = 8'h01;
Memory[4280] = 8'h13;
Memory[4287] = 8'h00;
Memory[4286] = 8'h0E;
Memory[4285] = 8'h8E;
Memory[4284] = 8'h13;
Memory[4291] = 8'h0D;
Memory[4290] = 8'h00;
Memory[4289] = 8'h10;
Memory[4288] = 8'h6F;
Memory[4295] = 8'h01;
Memory[4294] = 8'hC0;
Memory[4293] = 8'h01;
Memory[4292] = 8'h13;
Memory[4299] = 8'h00;
Memory[4298] = 8'h0E;
Memory[4297] = 8'h8E;
Memory[4296] = 8'h13;
Memory[4303] = 8'h7D;
Memory[4302] = 8'h50;
Memory[4301] = 8'h00;
Memory[4300] = 8'h6F;
Memory[4307] = 8'h01;
Memory[4306] = 8'hE0;
Memory[4305] = 8'h01;
Memory[4304] = 8'h13;
Memory[4311] = 8'h19;
Memory[4310] = 8'h0B;
Memory[4309] = 8'h21;
Memory[4308] = 8'h83;
Memory[4315] = 8'h19;
Memory[4314] = 8'h4B;
Memory[4313] = 8'h22;
Memory[4312] = 8'h03;
Memory[4319] = 8'h00;
Memory[4318] = 8'h00;
Memory[4317] = 8'h02;
Memory[4316] = 8'h93;
Memory[4323] = 8'hFF;
Memory[4322] = 8'hF0;
Memory[4321] = 8'h03;
Memory[4320] = 8'h13;
Memory[4327] = 8'h00;
Memory[4326] = 8'h83;
Memory[4325] = 8'h53;
Memory[4324] = 8'h13;
Memory[4331] = 8'h00;
Memory[4330] = 8'h3B;
Memory[4329] = 8'h20;
Memory[4328] = 8'h23;
Memory[4335] = 8'h00;
Memory[4334] = 8'h4B;
Memory[4333] = 8'h22;
Memory[4332] = 8'h23;
Memory[4339] = 8'h01;
Memory[4338] = 8'hDE;
Memory[4337] = 8'h14;
Memory[4336] = 8'h63;
Memory[4343] = 8'h09;
Memory[4342] = 8'hC0;
Memory[4341] = 8'h00;
Memory[4340] = 8'h6F;
Memory[4347] = 8'h01;
Memory[4346] = 8'hDE;
Memory[4345] = 8'h42;
Memory[4344] = 8'h33;
Memory[4351] = 8'h01;
Memory[4350] = 8'h82;
Memory[4349] = 8'h71;
Memory[4348] = 8'hB3;
Memory[4355] = 8'h01;
Memory[4354] = 8'hD1;
Memory[4353] = 8'hF1;
Memory[4352] = 8'hB3;
Memory[4359] = 8'h00;
Memory[4358] = 8'h01;
Memory[4357] = 8'h84;
Memory[4356] = 8'h63;
Memory[4363] = 8'h0D;
Memory[4362] = 8'h00;
Memory[4361] = 8'h20;
Memory[4360] = 8'h6F;
Memory[4367] = 8'hFF;
Memory[4366] = 8'hF2;
Memory[4365] = 8'h71;
Memory[4364] = 8'h93;
Memory[4371] = 8'h01;
Memory[4370] = 8'hD1;
Memory[4369] = 8'hF1;
Memory[4368] = 8'hB3;
Memory[4375] = 8'h00;
Memory[4374] = 8'h01;
Memory[4373] = 8'h94;
Memory[4372] = 8'h63;
Memory[4379] = 8'h2C;
Memory[4378] = 8'h40;
Memory[4377] = 8'h00;
Memory[4376] = 8'h6F;
Memory[4383] = 8'h40;
Memory[4382] = 8'h00;
Memory[4381] = 8'h02;
Memory[4380] = 8'h13;
Memory[4387] = 8'h00;
Memory[4386] = 8'h12;
Memory[4385] = 8'h12;
Memory[4384] = 8'h13;
Memory[4391] = 8'h00;
Memory[4390] = 8'h41;
Memory[4389] = 8'hF2;
Memory[4388] = 8'h33;
Memory[4395] = 8'h08;
Memory[4394] = 8'h02;
Memory[4393] = 8'h10;
Memory[4392] = 8'h63;
Memory[4399] = 8'h40;
Memory[4398] = 8'h01;
Memory[4397] = 8'hF2;
Memory[4396] = 8'h13;
Memory[4403] = 8'h08;
Memory[4402] = 8'h02;
Memory[4401] = 8'h1C;
Memory[4400] = 8'h63;
Memory[4407] = 8'h20;
Memory[4406] = 8'h01;
Memory[4405] = 8'hF2;
Memory[4404] = 8'h13;
Memory[4411] = 8'h0A;
Memory[4410] = 8'h02;
Memory[4409] = 8'h18;
Memory[4408] = 8'h63;
Memory[4415] = 8'h10;
Memory[4414] = 8'h01;
Memory[4413] = 8'hF2;
Memory[4412] = 8'h13;
Memory[4419] = 8'h0C;
Memory[4418] = 8'h02;
Memory[4417] = 8'h14;
Memory[4416] = 8'h63;
Memory[4423] = 8'h08;
Memory[4422] = 8'h01;
Memory[4421] = 8'hF2;
Memory[4420] = 8'h13;
Memory[4427] = 8'h0E;
Memory[4426] = 8'h02;
Memory[4425] = 8'h10;
Memory[4424] = 8'h63;
Memory[4431] = 8'h04;
Memory[4430] = 8'h01;
Memory[4429] = 8'hF2;
Memory[4428] = 8'h13;
Memory[4435] = 8'h0E;
Memory[4434] = 8'h02;
Memory[4433] = 8'h1C;
Memory[4432] = 8'h63;
Memory[4439] = 8'h02;
Memory[4438] = 8'h01;
Memory[4437] = 8'hF2;
Memory[4436] = 8'h13;
Memory[4443] = 8'h10;
Memory[4442] = 8'h02;
Memory[4441] = 8'h18;
Memory[4440] = 8'h63;
Memory[4447] = 8'h01;
Memory[4446] = 8'h01;
Memory[4445] = 8'hF2;
Memory[4444] = 8'h13;
Memory[4451] = 8'h12;
Memory[4450] = 8'h02;
Memory[4449] = 8'h14;
Memory[4448] = 8'h63;
Memory[4455] = 8'h00;
Memory[4454] = 8'h81;
Memory[4453] = 8'hF2;
Memory[4452] = 8'h13;
Memory[4459] = 8'h14;
Memory[4458] = 8'h02;
Memory[4457] = 8'h10;
Memory[4456] = 8'h63;
Memory[4463] = 8'h00;
Memory[4462] = 8'h41;
Memory[4461] = 8'hF2;
Memory[4460] = 8'h13;
Memory[4467] = 8'h14;
Memory[4466] = 8'h02;
Memory[4465] = 8'h1C;
Memory[4464] = 8'h63;
Memory[4471] = 8'h00;
Memory[4470] = 8'h21;
Memory[4469] = 8'hF2;
Memory[4468] = 8'h13;
Memory[4475] = 8'h00;
Memory[4474] = 8'h02;
Memory[4473] = 8'h18;
Memory[4472] = 8'h63;
Memory[4479] = 8'h00;
Memory[4478] = 8'h11;
Memory[4477] = 8'hF2;
Memory[4476] = 8'h13;
Memory[4483] = 8'h18;
Memory[4482] = 8'h02;
Memory[4481] = 8'h1C;
Memory[4480] = 8'h63;
Memory[4487] = 8'h2C;
Memory[4486] = 8'h40;
Memory[4485] = 8'h00;
Memory[4484] = 8'h6F;
Memory[4491] = 8'h00;
Memory[4490] = 8'h82;
Memory[4489] = 8'h92;
Memory[4488] = 8'h93;
Memory[4495] = 8'h00;
Memory[4494] = 8'h02;
Memory[4493] = 8'h82;
Memory[4492] = 8'h93;
Memory[4499] = 8'h00;
Memory[4498] = 8'h62;
Memory[4497] = 8'hF2;
Memory[4496] = 8'hB3;
Memory[4503] = 8'h19;
Memory[4502] = 8'h4B;
Memory[4501] = 8'h22;
Memory[4500] = 8'h03;
Memory[4507] = 8'h00;
Memory[4506] = 8'h52;
Memory[4505] = 8'h02;
Memory[4504] = 8'h33;
Memory[4511] = 8'h00;
Memory[4510] = 8'h4B;
Memory[4509] = 8'h22;
Memory[4508] = 8'h23;
Memory[4515] = 8'h00;
Memory[4514] = 8'h0E;
Memory[4513] = 8'h8E;
Memory[4512] = 8'h13;
Memory[4519] = 8'h2C;
Memory[4518] = 8'h40;
Memory[4517] = 8'h00;
Memory[4516] = 8'h6F;
Memory[4523] = 8'h00;
Memory[4522] = 8'h82;
Memory[4521] = 8'h92;
Memory[4520] = 8'h93;
Memory[4527] = 8'h00;
Memory[4526] = 8'h12;
Memory[4525] = 8'h82;
Memory[4524] = 8'h93;
Memory[4531] = 8'h00;
Memory[4530] = 8'h62;
Memory[4529] = 8'hF2;
Memory[4528] = 8'hB3;
Memory[4535] = 8'h19;
Memory[4534] = 8'h4B;
Memory[4533] = 8'h22;
Memory[4532] = 8'h03;
Memory[4539] = 8'h00;
Memory[4538] = 8'h52;
Memory[4537] = 8'h02;
Memory[4536] = 8'h33;
Memory[4543] = 8'h00;
Memory[4542] = 8'h4B;
Memory[4541] = 8'h22;
Memory[4540] = 8'h23;
Memory[4547] = 8'h00;
Memory[4546] = 8'h0E;
Memory[4545] = 8'h8E;
Memory[4544] = 8'h13;
Memory[4551] = 8'h2C;
Memory[4550] = 8'h40;
Memory[4549] = 8'h00;
Memory[4548] = 8'h6F;
Memory[4555] = 8'h00;
Memory[4554] = 8'h82;
Memory[4553] = 8'h92;
Memory[4552] = 8'h93;
Memory[4559] = 8'h00;
Memory[4558] = 8'h22;
Memory[4557] = 8'h82;
Memory[4556] = 8'h93;
Memory[4563] = 8'h00;
Memory[4562] = 8'h62;
Memory[4561] = 8'hF2;
Memory[4560] = 8'hB3;
Memory[4567] = 8'h19;
Memory[4566] = 8'h4B;
Memory[4565] = 8'h22;
Memory[4564] = 8'h03;
Memory[4571] = 8'h00;
Memory[4570] = 8'h52;
Memory[4569] = 8'h02;
Memory[4568] = 8'h33;
Memory[4575] = 8'h00;
Memory[4574] = 8'h4B;
Memory[4573] = 8'h22;
Memory[4572] = 8'h23;
Memory[4579] = 8'h00;
Memory[4578] = 8'h0E;
Memory[4577] = 8'h8E;
Memory[4576] = 8'h13;
Memory[4583] = 8'h2C;
Memory[4582] = 8'h40;
Memory[4581] = 8'h00;
Memory[4580] = 8'h6F;
Memory[4587] = 8'h00;
Memory[4586] = 8'h82;
Memory[4585] = 8'h92;
Memory[4584] = 8'h93;
Memory[4591] = 8'h00;
Memory[4590] = 8'h32;
Memory[4589] = 8'h82;
Memory[4588] = 8'h93;
Memory[4595] = 8'h00;
Memory[4594] = 8'h62;
Memory[4593] = 8'hF2;
Memory[4592] = 8'hB3;
Memory[4599] = 8'h19;
Memory[4598] = 8'h4B;
Memory[4597] = 8'h22;
Memory[4596] = 8'h03;
Memory[4603] = 8'h00;
Memory[4602] = 8'h52;
Memory[4601] = 8'h02;
Memory[4600] = 8'h33;
Memory[4607] = 8'h00;
Memory[4606] = 8'h4B;
Memory[4605] = 8'h22;
Memory[4604] = 8'h23;
Memory[4611] = 8'h00;
Memory[4610] = 8'h0E;
Memory[4609] = 8'h8E;
Memory[4608] = 8'h13;
Memory[4615] = 8'h2C;
Memory[4614] = 8'h40;
Memory[4613] = 8'h00;
Memory[4612] = 8'h6F;
Memory[4619] = 8'h00;
Memory[4618] = 8'h82;
Memory[4617] = 8'h92;
Memory[4616] = 8'h93;
Memory[4623] = 8'h00;
Memory[4622] = 8'h42;
Memory[4621] = 8'h82;
Memory[4620] = 8'h93;
Memory[4627] = 8'h00;
Memory[4626] = 8'h62;
Memory[4625] = 8'hF2;
Memory[4624] = 8'hB3;
Memory[4631] = 8'h19;
Memory[4630] = 8'h4B;
Memory[4629] = 8'h22;
Memory[4628] = 8'h03;
Memory[4635] = 8'h00;
Memory[4634] = 8'h52;
Memory[4633] = 8'h02;
Memory[4632] = 8'h33;
Memory[4639] = 8'h00;
Memory[4638] = 8'h4B;
Memory[4637] = 8'h22;
Memory[4636] = 8'h23;
Memory[4643] = 8'h00;
Memory[4642] = 8'h0E;
Memory[4641] = 8'h8E;
Memory[4640] = 8'h13;
Memory[4647] = 8'h2C;
Memory[4646] = 8'h40;
Memory[4645] = 8'h00;
Memory[4644] = 8'h6F;
Memory[4651] = 8'h00;
Memory[4650] = 8'h82;
Memory[4649] = 8'h92;
Memory[4648] = 8'h93;
Memory[4655] = 8'h00;
Memory[4654] = 8'h52;
Memory[4653] = 8'h82;
Memory[4652] = 8'h93;
Memory[4659] = 8'h00;
Memory[4658] = 8'h62;
Memory[4657] = 8'hF2;
Memory[4656] = 8'hB3;
Memory[4663] = 8'h19;
Memory[4662] = 8'h4B;
Memory[4661] = 8'h22;
Memory[4660] = 8'h03;
Memory[4667] = 8'h00;
Memory[4666] = 8'h52;
Memory[4665] = 8'h02;
Memory[4664] = 8'h33;
Memory[4671] = 8'h00;
Memory[4670] = 8'h4B;
Memory[4669] = 8'h22;
Memory[4668] = 8'h23;
Memory[4675] = 8'h00;
Memory[4674] = 8'h0E;
Memory[4673] = 8'h8E;
Memory[4672] = 8'h13;
Memory[4679] = 8'h2C;
Memory[4678] = 8'h40;
Memory[4677] = 8'h00;
Memory[4676] = 8'h6F;
Memory[4683] = 8'h00;
Memory[4682] = 8'h82;
Memory[4681] = 8'h92;
Memory[4680] = 8'h93;
Memory[4687] = 8'h00;
Memory[4686] = 8'h62;
Memory[4685] = 8'h82;
Memory[4684] = 8'h93;
Memory[4691] = 8'h00;
Memory[4690] = 8'h62;
Memory[4689] = 8'hF2;
Memory[4688] = 8'hB3;
Memory[4695] = 8'h19;
Memory[4694] = 8'h4B;
Memory[4693] = 8'h22;
Memory[4692] = 8'h03;
Memory[4699] = 8'h00;
Memory[4698] = 8'h52;
Memory[4697] = 8'h02;
Memory[4696] = 8'h33;
Memory[4703] = 8'h00;
Memory[4702] = 8'h4B;
Memory[4701] = 8'h22;
Memory[4700] = 8'h23;
Memory[4707] = 8'h00;
Memory[4706] = 8'h0E;
Memory[4705] = 8'h8E;
Memory[4704] = 8'h13;
Memory[4711] = 8'h2C;
Memory[4710] = 8'h40;
Memory[4709] = 8'h00;
Memory[4708] = 8'h6F;
Memory[4715] = 8'h00;
Memory[4714] = 8'h82;
Memory[4713] = 8'h92;
Memory[4712] = 8'h93;
Memory[4719] = 8'h00;
Memory[4718] = 8'h72;
Memory[4717] = 8'h82;
Memory[4716] = 8'h93;
Memory[4723] = 8'h00;
Memory[4722] = 8'h62;
Memory[4721] = 8'hF2;
Memory[4720] = 8'hB3;
Memory[4727] = 8'h19;
Memory[4726] = 8'h4B;
Memory[4725] = 8'h22;
Memory[4724] = 8'h03;
Memory[4731] = 8'h00;
Memory[4730] = 8'h52;
Memory[4729] = 8'h02;
Memory[4728] = 8'h33;
Memory[4735] = 8'h00;
Memory[4734] = 8'h4B;
Memory[4733] = 8'h22;
Memory[4732] = 8'h23;
Memory[4739] = 8'h00;
Memory[4738] = 8'h0E;
Memory[4737] = 8'h8E;
Memory[4736] = 8'h13;
Memory[4743] = 8'h2C;
Memory[4742] = 8'h40;
Memory[4741] = 8'h00;
Memory[4740] = 8'h6F;
Memory[4747] = 8'h00;
Memory[4746] = 8'h82;
Memory[4745] = 8'h92;
Memory[4744] = 8'h93;
Memory[4751] = 8'h00;
Memory[4750] = 8'h82;
Memory[4749] = 8'h82;
Memory[4748] = 8'h93;
Memory[4755] = 8'h00;
Memory[4754] = 8'h62;
Memory[4753] = 8'hF2;
Memory[4752] = 8'hB3;
Memory[4759] = 8'h19;
Memory[4758] = 8'h4B;
Memory[4757] = 8'h22;
Memory[4756] = 8'h03;
Memory[4763] = 8'h00;
Memory[4762] = 8'h52;
Memory[4761] = 8'h02;
Memory[4760] = 8'h33;
Memory[4767] = 8'h00;
Memory[4766] = 8'h4B;
Memory[4765] = 8'h22;
Memory[4764] = 8'h23;
Memory[4771] = 8'h00;
Memory[4770] = 8'h0E;
Memory[4769] = 8'h8E;
Memory[4768] = 8'h13;
Memory[4775] = 8'h2C;
Memory[4774] = 8'h40;
Memory[4773] = 8'h00;
Memory[4772] = 8'h6F;
Memory[4779] = 8'h00;
Memory[4778] = 8'h82;
Memory[4777] = 8'h92;
Memory[4776] = 8'h93;
Memory[4783] = 8'h00;
Memory[4782] = 8'h92;
Memory[4781] = 8'h82;
Memory[4780] = 8'h93;
Memory[4787] = 8'h00;
Memory[4786] = 8'h62;
Memory[4785] = 8'hF2;
Memory[4784] = 8'hB3;
Memory[4791] = 8'h19;
Memory[4790] = 8'h4B;
Memory[4789] = 8'h22;
Memory[4788] = 8'h03;
Memory[4795] = 8'h00;
Memory[4794] = 8'h52;
Memory[4793] = 8'h02;
Memory[4792] = 8'h33;
Memory[4799] = 8'h00;
Memory[4798] = 8'h4B;
Memory[4797] = 8'h22;
Memory[4796] = 8'h23;
Memory[4803] = 8'h00;
Memory[4802] = 8'h0E;
Memory[4801] = 8'h8E;
Memory[4800] = 8'h13;
Memory[4807] = 8'h2C;
Memory[4806] = 8'h40;
Memory[4805] = 8'h00;
Memory[4804] = 8'h6F;
Memory[4811] = 8'h01;
Memory[4810] = 8'hD0;
Memory[4809] = 8'h01;
Memory[4808] = 8'h13;
Memory[4815] = 8'h00;
Memory[4814] = 8'h0E;
Memory[4813] = 8'h8E;
Memory[4812] = 8'h13;
Memory[4819] = 8'h0F;
Memory[4818] = 8'hF0;
Memory[4817] = 8'h01;
Memory[4816] = 8'h93;
Memory[4823] = 8'h01;
Memory[4822] = 8'h01;
Memory[4821] = 8'h91;
Memory[4820] = 8'h93;
Memory[4827] = 8'h00;
Memory[4826] = 8'h32;
Memory[4825] = 8'hF1;
Memory[4824] = 8'hB3;
Memory[4831] = 8'h01;
Memory[4830] = 8'h01;
Memory[4829] = 8'hD1;
Memory[4828] = 8'h93;
Memory[4835] = 8'h06;
Memory[4834] = 8'h40;
Memory[4833] = 8'h02;
Memory[4832] = 8'h13;
Memory[4839] = 8'h02;
Memory[4838] = 8'h41;
Memory[4837] = 8'h82;
Memory[4836] = 8'h33;
Memory[4843] = 8'h0F;
Memory[4842] = 8'hF0;
Memory[4841] = 8'h01;
Memory[4840] = 8'h93;
Memory[4847] = 8'h00;
Memory[4846] = 8'h81;
Memory[4845] = 8'h91;
Memory[4844] = 8'h93;
Memory[4851] = 8'h00;
Memory[4850] = 8'h32;
Memory[4849] = 8'hF1;
Memory[4848] = 8'hB3;
Memory[4855] = 8'h00;
Memory[4854] = 8'h81;
Memory[4853] = 8'hD1;
Memory[4852] = 8'h93;
Memory[4859] = 8'h00;
Memory[4858] = 8'hA0;
Memory[4857] = 8'h03;
Memory[4856] = 8'h13;
Memory[4863] = 8'h02;
Memory[4862] = 8'h61;
Memory[4861] = 8'h81;
Memory[4860] = 8'hB3;
Memory[4867] = 8'h00;
Memory[4866] = 8'h41;
Memory[4865] = 8'h82;
Memory[4864] = 8'h33;
Memory[4871] = 8'h0F;
Memory[4870] = 8'hF0;
Memory[4869] = 8'h01;
Memory[4868] = 8'h93;
Memory[4875] = 8'h00;
Memory[4874] = 8'h32;
Memory[4873] = 8'hF1;
Memory[4872] = 8'hB3;
Memory[4879] = 8'h00;
Memory[4878] = 8'h41;
Memory[4877] = 8'h81;
Memory[4876] = 8'hB3;
Memory[4883] = 8'h00;
Memory[4882] = 8'h3B;
Memory[4881] = 8'h2C;
Memory[4880] = 8'h23;
Memory[4887] = 8'h04;
Memory[4886] = 8'h80;
Memory[4885] = 8'h10;
Memory[4884] = 8'h6F;
Memory[4891] = 8'h01;
Memory[4890] = 8'hD0;
Memory[4889] = 8'h01;
Memory[4888] = 8'h13;
Memory[4895] = 8'h00;
Memory[4894] = 8'h0E;
Memory[4893] = 8'h8E;
Memory[4892] = 8'h13;
Memory[4899] = 8'h04;
Memory[4898] = 8'h80;
Memory[4897] = 8'h10;
Memory[4896] = 8'h6F;
Memory[4903] = 8'h01;
Memory[4902] = 8'hF0;
Memory[4901] = 8'h01;
Memory[4900] = 8'h13;
Memory[4907] = 8'h19;
Memory[4906] = 8'h8B;
Memory[4905] = 8'h21;
Memory[4904] = 8'h83;
Memory[4911] = 8'h19;
Memory[4910] = 8'hCB;
Memory[4909] = 8'h22;
Memory[4908] = 8'h03;
Memory[4915] = 8'h01;
Memory[4914] = 8'hA0;
Memory[4913] = 8'h02;
Memory[4912] = 8'h93;
Memory[4919] = 8'h00;
Memory[4918] = 8'h3B;
Memory[4917] = 8'h20;
Memory[4916] = 8'h23;
Memory[4923] = 8'h00;
Memory[4922] = 8'h4B;
Memory[4921] = 8'h22;
Memory[4920] = 8'h23;
Memory[4927] = 8'h00;
Memory[4926] = 8'h5B;
Memory[4925] = 8'h24;
Memory[4924] = 8'h23;
Memory[4931] = 8'h01;
Memory[4930] = 8'hDE;
Memory[4929] = 8'h14;
Memory[4928] = 8'h63;
Memory[4935] = 8'h09;
Memory[4934] = 8'hC0;
Memory[4933] = 8'h00;
Memory[4932] = 8'h6F;
Memory[4939] = 8'h01;
Memory[4938] = 8'hDE;
Memory[4937] = 8'h42;
Memory[4936] = 8'h33;
Memory[4943] = 8'h01;
Memory[4942] = 8'h82;
Memory[4941] = 8'h71;
Memory[4940] = 8'hB3;
Memory[4947] = 8'h01;
Memory[4946] = 8'hD1;
Memory[4945] = 8'hF1;
Memory[4944] = 8'hB3;
Memory[4951] = 8'h00;
Memory[4950] = 8'h01;
Memory[4949] = 8'h84;
Memory[4948] = 8'h63;
Memory[4955] = 8'h0D;
Memory[4954] = 8'h00;
Memory[4953] = 8'h20;
Memory[4952] = 8'h6F;
Memory[4959] = 8'hFF;
Memory[4958] = 8'hF2;
Memory[4957] = 8'h71;
Memory[4956] = 8'h93;
Memory[4963] = 8'h01;
Memory[4962] = 8'hD1;
Memory[4961] = 8'hF1;
Memory[4960] = 8'hB3;
Memory[4967] = 8'h00;
Memory[4966] = 8'h01;
Memory[4965] = 8'h94;
Memory[4964] = 8'h63;
Memory[4971] = 8'h2C;
Memory[4970] = 8'h40;
Memory[4969] = 8'h00;
Memory[4968] = 8'h6F;
Memory[4975] = 8'h40;
Memory[4974] = 8'h01;
Memory[4973] = 8'hF2;
Memory[4972] = 8'h13;
Memory[4979] = 8'h00;
Memory[4978] = 8'h02;
Memory[4977] = 8'h1C;
Memory[4976] = 8'h63;
Memory[4983] = 8'h00;
Memory[4982] = 8'h41;
Memory[4981] = 8'hF2;
Memory[4980] = 8'h13;
Memory[4987] = 8'h00;
Memory[4986] = 8'h02;
Memory[4985] = 8'h1E;
Memory[4984] = 8'h63;
Memory[4991] = 8'h00;
Memory[4990] = 8'h11;
Memory[4989] = 8'hF2;
Memory[4988] = 8'h13;
Memory[4995] = 8'h02;
Memory[4994] = 8'h02;
Memory[4993] = 8'h10;
Memory[4992] = 8'h63;
Memory[4999] = 8'h2C;
Memory[4998] = 8'h40;
Memory[4997] = 8'h00;
Memory[4996] = 8'h6F;
Memory[5003] = 8'h01;
Memory[5002] = 8'hD0;
Memory[5001] = 8'h01;
Memory[5000] = 8'h13;
Memory[5007] = 8'h00;
Memory[5006] = 8'h0E;
Memory[5005] = 8'h8E;
Memory[5004] = 8'h13;
Memory[5011] = 8'h04;
Memory[5010] = 8'h80;
Memory[5009] = 8'h10;
Memory[5008] = 8'h6F;
Memory[5015] = 8'h02;
Memory[5014] = 8'h00;
Memory[5013] = 8'h01;
Memory[5012] = 8'h13;
Memory[5019] = 8'h00;
Memory[5018] = 8'h0E;
Memory[5017] = 8'h8E;
Memory[5016] = 8'h13;
Memory[5023] = 8'h3A;
Memory[5022] = 8'hC0;
Memory[5021] = 8'h10;
Memory[5020] = 8'h6F;
Memory[5027] = 8'h02;
Memory[5026] = 8'h10;
Memory[5025] = 8'h01;
Memory[5024] = 8'h13;
Memory[5031] = 8'h00;
Memory[5030] = 8'h0E;
Memory[5029] = 8'h8E;
Memory[5028] = 8'h13;
Memory[5035] = 8'h60;
Memory[5034] = 8'h00;
Memory[5033] = 8'h10;
Memory[5032] = 8'h6F;
Memory[5039] = 8'h02;
Memory[5038] = 8'h00;
Memory[5037] = 8'h01;
Memory[5036] = 8'h13;
Memory[5043] = 8'h25;
Memory[5042] = 8'h8B;
Memory[5041] = 8'h21;
Memory[5040] = 8'h83;
Memory[5047] = 8'h25;
Memory[5046] = 8'hCB;
Memory[5045] = 8'h22;
Memory[5044] = 8'h03;
Memory[5051] = 8'h00;
Memory[5050] = 8'h00;
Memory[5049] = 8'h02;
Memory[5048] = 8'h93;
Memory[5055] = 8'hFF;
Memory[5054] = 8'hF0;
Memory[5053] = 8'h03;
Memory[5052] = 8'h13;
Memory[5059] = 8'h00;
Memory[5058] = 8'h83;
Memory[5057] = 8'h53;
Memory[5056] = 8'h13;
Memory[5063] = 8'h00;
Memory[5062] = 8'h3B;
Memory[5061] = 8'h20;
Memory[5060] = 8'h23;
Memory[5067] = 8'h00;
Memory[5066] = 8'h4B;
Memory[5065] = 8'h22;
Memory[5064] = 8'h23;
Memory[5071] = 8'h01;
Memory[5070] = 8'hDE;
Memory[5069] = 8'h14;
Memory[5068] = 8'h63;
Memory[5075] = 8'h09;
Memory[5074] = 8'hC0;
Memory[5073] = 8'h00;
Memory[5072] = 8'h6F;
Memory[5079] = 8'h01;
Memory[5078] = 8'hDE;
Memory[5077] = 8'h42;
Memory[5076] = 8'h33;
Memory[5083] = 8'h01;
Memory[5082] = 8'h82;
Memory[5081] = 8'h71;
Memory[5080] = 8'hB3;
Memory[5087] = 8'h01;
Memory[5086] = 8'hD1;
Memory[5085] = 8'hF1;
Memory[5084] = 8'hB3;
Memory[5091] = 8'h00;
Memory[5090] = 8'h01;
Memory[5089] = 8'h84;
Memory[5088] = 8'h63;
Memory[5095] = 8'h0D;
Memory[5094] = 8'h00;
Memory[5093] = 8'h20;
Memory[5092] = 8'h6F;
Memory[5099] = 8'hFF;
Memory[5098] = 8'hF2;
Memory[5097] = 8'h71;
Memory[5096] = 8'h93;
Memory[5103] = 8'h01;
Memory[5102] = 8'hD1;
Memory[5101] = 8'hF1;
Memory[5100] = 8'hB3;
Memory[5107] = 8'h00;
Memory[5106] = 8'h01;
Memory[5105] = 8'h94;
Memory[5104] = 8'h63;
Memory[5111] = 8'h2C;
Memory[5110] = 8'h40;
Memory[5109] = 8'h00;
Memory[5108] = 8'h6F;
Memory[5115] = 8'h40;
Memory[5114] = 8'h00;
Memory[5113] = 8'h02;
Memory[5112] = 8'h13;
Memory[5119] = 8'h00;
Memory[5118] = 8'h12;
Memory[5117] = 8'h12;
Memory[5116] = 8'h13;
Memory[5123] = 8'h00;
Memory[5122] = 8'h41;
Memory[5121] = 8'hF2;
Memory[5120] = 8'h33;
Memory[5127] = 8'h08;
Memory[5126] = 8'h02;
Memory[5125] = 8'h10;
Memory[5124] = 8'h63;
Memory[5131] = 8'h40;
Memory[5130] = 8'h01;
Memory[5129] = 8'hF2;
Memory[5128] = 8'h13;
Memory[5135] = 8'h08;
Memory[5134] = 8'h02;
Memory[5133] = 8'h1C;
Memory[5132] = 8'h63;
Memory[5139] = 8'h20;
Memory[5138] = 8'h01;
Memory[5137] = 8'hF2;
Memory[5136] = 8'h13;
Memory[5143] = 8'h0A;
Memory[5142] = 8'h02;
Memory[5141] = 8'h18;
Memory[5140] = 8'h63;
Memory[5147] = 8'h10;
Memory[5146] = 8'h01;
Memory[5145] = 8'hF2;
Memory[5144] = 8'h13;
Memory[5151] = 8'h0C;
Memory[5150] = 8'h02;
Memory[5149] = 8'h14;
Memory[5148] = 8'h63;
Memory[5155] = 8'h08;
Memory[5154] = 8'h01;
Memory[5153] = 8'hF2;
Memory[5152] = 8'h13;
Memory[5159] = 8'h0E;
Memory[5158] = 8'h02;
Memory[5157] = 8'h10;
Memory[5156] = 8'h63;
Memory[5163] = 8'h04;
Memory[5162] = 8'h01;
Memory[5161] = 8'hF2;
Memory[5160] = 8'h13;
Memory[5167] = 8'h0E;
Memory[5166] = 8'h02;
Memory[5165] = 8'h1C;
Memory[5164] = 8'h63;
Memory[5171] = 8'h02;
Memory[5170] = 8'h01;
Memory[5169] = 8'hF2;
Memory[5168] = 8'h13;
Memory[5175] = 8'h10;
Memory[5174] = 8'h02;
Memory[5173] = 8'h18;
Memory[5172] = 8'h63;
Memory[5179] = 8'h01;
Memory[5178] = 8'h01;
Memory[5177] = 8'hF2;
Memory[5176] = 8'h13;
Memory[5183] = 8'h12;
Memory[5182] = 8'h02;
Memory[5181] = 8'h14;
Memory[5180] = 8'h63;
Memory[5187] = 8'h00;
Memory[5186] = 8'h81;
Memory[5185] = 8'hF2;
Memory[5184] = 8'h13;
Memory[5191] = 8'h14;
Memory[5190] = 8'h02;
Memory[5189] = 8'h10;
Memory[5188] = 8'h63;
Memory[5195] = 8'h00;
Memory[5194] = 8'h41;
Memory[5193] = 8'hF2;
Memory[5192] = 8'h13;
Memory[5199] = 8'h14;
Memory[5198] = 8'h02;
Memory[5197] = 8'h1C;
Memory[5196] = 8'h63;
Memory[5203] = 8'h00;
Memory[5202] = 8'h21;
Memory[5201] = 8'hF2;
Memory[5200] = 8'h13;
Memory[5207] = 8'h00;
Memory[5206] = 8'h02;
Memory[5205] = 8'h18;
Memory[5204] = 8'h63;
Memory[5211] = 8'h00;
Memory[5210] = 8'h11;
Memory[5209] = 8'hF2;
Memory[5208] = 8'h13;
Memory[5215] = 8'h18;
Memory[5214] = 8'h02;
Memory[5213] = 8'h1C;
Memory[5212] = 8'h63;
Memory[5219] = 8'h2C;
Memory[5218] = 8'h40;
Memory[5217] = 8'h00;
Memory[5216] = 8'h6F;
Memory[5223] = 8'h00;
Memory[5222] = 8'h82;
Memory[5221] = 8'h92;
Memory[5220] = 8'h93;
Memory[5227] = 8'h00;
Memory[5226] = 8'h02;
Memory[5225] = 8'h82;
Memory[5224] = 8'h93;
Memory[5231] = 8'h00;
Memory[5230] = 8'h62;
Memory[5229] = 8'hF2;
Memory[5228] = 8'hB3;
Memory[5235] = 8'h25;
Memory[5234] = 8'hCB;
Memory[5233] = 8'h22;
Memory[5232] = 8'h03;
Memory[5239] = 8'h00;
Memory[5238] = 8'h52;
Memory[5237] = 8'h02;
Memory[5236] = 8'h33;
Memory[5243] = 8'h00;
Memory[5242] = 8'h4B;
Memory[5241] = 8'h22;
Memory[5240] = 8'h23;
Memory[5247] = 8'h00;
Memory[5246] = 8'h0E;
Memory[5245] = 8'h8E;
Memory[5244] = 8'h13;
Memory[5251] = 8'h2C;
Memory[5250] = 8'h40;
Memory[5249] = 8'h00;
Memory[5248] = 8'h6F;
Memory[5255] = 8'h00;
Memory[5254] = 8'h82;
Memory[5253] = 8'h92;
Memory[5252] = 8'h93;
Memory[5259] = 8'h00;
Memory[5258] = 8'h12;
Memory[5257] = 8'h82;
Memory[5256] = 8'h93;
Memory[5263] = 8'h00;
Memory[5262] = 8'h62;
Memory[5261] = 8'hF2;
Memory[5260] = 8'hB3;
Memory[5267] = 8'h25;
Memory[5266] = 8'hCB;
Memory[5265] = 8'h22;
Memory[5264] = 8'h03;
Memory[5271] = 8'h00;
Memory[5270] = 8'h52;
Memory[5269] = 8'h02;
Memory[5268] = 8'h33;
Memory[5275] = 8'h00;
Memory[5274] = 8'h4B;
Memory[5273] = 8'h22;
Memory[5272] = 8'h23;
Memory[5279] = 8'h00;
Memory[5278] = 8'h0E;
Memory[5277] = 8'h8E;
Memory[5276] = 8'h13;
Memory[5283] = 8'h2C;
Memory[5282] = 8'h40;
Memory[5281] = 8'h00;
Memory[5280] = 8'h6F;
Memory[5287] = 8'h00;
Memory[5286] = 8'h82;
Memory[5285] = 8'h92;
Memory[5284] = 8'h93;
Memory[5291] = 8'h00;
Memory[5290] = 8'h22;
Memory[5289] = 8'h82;
Memory[5288] = 8'h93;
Memory[5295] = 8'h00;
Memory[5294] = 8'h62;
Memory[5293] = 8'hF2;
Memory[5292] = 8'hB3;
Memory[5299] = 8'h25;
Memory[5298] = 8'hCB;
Memory[5297] = 8'h22;
Memory[5296] = 8'h03;
Memory[5303] = 8'h00;
Memory[5302] = 8'h52;
Memory[5301] = 8'h02;
Memory[5300] = 8'h33;
Memory[5307] = 8'h00;
Memory[5306] = 8'h4B;
Memory[5305] = 8'h22;
Memory[5304] = 8'h23;
Memory[5311] = 8'h00;
Memory[5310] = 8'h0E;
Memory[5309] = 8'h8E;
Memory[5308] = 8'h13;
Memory[5315] = 8'h2C;
Memory[5314] = 8'h40;
Memory[5313] = 8'h00;
Memory[5312] = 8'h6F;
Memory[5319] = 8'h00;
Memory[5318] = 8'h82;
Memory[5317] = 8'h92;
Memory[5316] = 8'h93;
Memory[5323] = 8'h00;
Memory[5322] = 8'h32;
Memory[5321] = 8'h82;
Memory[5320] = 8'h93;
Memory[5327] = 8'h00;
Memory[5326] = 8'h62;
Memory[5325] = 8'hF2;
Memory[5324] = 8'hB3;
Memory[5331] = 8'h25;
Memory[5330] = 8'hCB;
Memory[5329] = 8'h22;
Memory[5328] = 8'h03;
Memory[5335] = 8'h00;
Memory[5334] = 8'h52;
Memory[5333] = 8'h02;
Memory[5332] = 8'h33;
Memory[5339] = 8'h00;
Memory[5338] = 8'h4B;
Memory[5337] = 8'h22;
Memory[5336] = 8'h23;
Memory[5343] = 8'h00;
Memory[5342] = 8'h0E;
Memory[5341] = 8'h8E;
Memory[5340] = 8'h13;
Memory[5347] = 8'h2C;
Memory[5346] = 8'h40;
Memory[5345] = 8'h00;
Memory[5344] = 8'h6F;
Memory[5351] = 8'h00;
Memory[5350] = 8'h82;
Memory[5349] = 8'h92;
Memory[5348] = 8'h93;
Memory[5355] = 8'h00;
Memory[5354] = 8'h42;
Memory[5353] = 8'h82;
Memory[5352] = 8'h93;
Memory[5359] = 8'h00;
Memory[5358] = 8'h62;
Memory[5357] = 8'hF2;
Memory[5356] = 8'hB3;
Memory[5363] = 8'h25;
Memory[5362] = 8'hCB;
Memory[5361] = 8'h22;
Memory[5360] = 8'h03;
Memory[5367] = 8'h00;
Memory[5366] = 8'h52;
Memory[5365] = 8'h02;
Memory[5364] = 8'h33;
Memory[5371] = 8'h00;
Memory[5370] = 8'h4B;
Memory[5369] = 8'h22;
Memory[5368] = 8'h23;
Memory[5375] = 8'h00;
Memory[5374] = 8'h0E;
Memory[5373] = 8'h8E;
Memory[5372] = 8'h13;
Memory[5379] = 8'h2C;
Memory[5378] = 8'h40;
Memory[5377] = 8'h00;
Memory[5376] = 8'h6F;
Memory[5383] = 8'h00;
Memory[5382] = 8'h82;
Memory[5381] = 8'h92;
Memory[5380] = 8'h93;
Memory[5387] = 8'h00;
Memory[5386] = 8'h52;
Memory[5385] = 8'h82;
Memory[5384] = 8'h93;
Memory[5391] = 8'h00;
Memory[5390] = 8'h62;
Memory[5389] = 8'hF2;
Memory[5388] = 8'hB3;
Memory[5395] = 8'h25;
Memory[5394] = 8'hCB;
Memory[5393] = 8'h22;
Memory[5392] = 8'h03;
Memory[5399] = 8'h00;
Memory[5398] = 8'h52;
Memory[5397] = 8'h02;
Memory[5396] = 8'h33;
Memory[5403] = 8'h00;
Memory[5402] = 8'h4B;
Memory[5401] = 8'h22;
Memory[5400] = 8'h23;
Memory[5407] = 8'h00;
Memory[5406] = 8'h0E;
Memory[5405] = 8'h8E;
Memory[5404] = 8'h13;
Memory[5411] = 8'h2C;
Memory[5410] = 8'h40;
Memory[5409] = 8'h00;
Memory[5408] = 8'h6F;
Memory[5415] = 8'h00;
Memory[5414] = 8'h82;
Memory[5413] = 8'h92;
Memory[5412] = 8'h93;
Memory[5419] = 8'h00;
Memory[5418] = 8'h62;
Memory[5417] = 8'h82;
Memory[5416] = 8'h93;
Memory[5423] = 8'h00;
Memory[5422] = 8'h62;
Memory[5421] = 8'hF2;
Memory[5420] = 8'hB3;
Memory[5427] = 8'h25;
Memory[5426] = 8'hCB;
Memory[5425] = 8'h22;
Memory[5424] = 8'h03;
Memory[5431] = 8'h00;
Memory[5430] = 8'h52;
Memory[5429] = 8'h02;
Memory[5428] = 8'h33;
Memory[5435] = 8'h00;
Memory[5434] = 8'h4B;
Memory[5433] = 8'h22;
Memory[5432] = 8'h23;
Memory[5439] = 8'h00;
Memory[5438] = 8'h0E;
Memory[5437] = 8'h8E;
Memory[5436] = 8'h13;
Memory[5443] = 8'h2C;
Memory[5442] = 8'h40;
Memory[5441] = 8'h00;
Memory[5440] = 8'h6F;
Memory[5447] = 8'h00;
Memory[5446] = 8'h82;
Memory[5445] = 8'h92;
Memory[5444] = 8'h93;
Memory[5451] = 8'h00;
Memory[5450] = 8'h72;
Memory[5449] = 8'h82;
Memory[5448] = 8'h93;
Memory[5455] = 8'h00;
Memory[5454] = 8'h62;
Memory[5453] = 8'hF2;
Memory[5452] = 8'hB3;
Memory[5459] = 8'h25;
Memory[5458] = 8'hCB;
Memory[5457] = 8'h22;
Memory[5456] = 8'h03;
Memory[5463] = 8'h00;
Memory[5462] = 8'h52;
Memory[5461] = 8'h02;
Memory[5460] = 8'h33;
Memory[5467] = 8'h00;
Memory[5466] = 8'h4B;
Memory[5465] = 8'h22;
Memory[5464] = 8'h23;
Memory[5471] = 8'h00;
Memory[5470] = 8'h0E;
Memory[5469] = 8'h8E;
Memory[5468] = 8'h13;
Memory[5475] = 8'h2C;
Memory[5474] = 8'h40;
Memory[5473] = 8'h00;
Memory[5472] = 8'h6F;
Memory[5479] = 8'h00;
Memory[5478] = 8'h82;
Memory[5477] = 8'h92;
Memory[5476] = 8'h93;
Memory[5483] = 8'h00;
Memory[5482] = 8'h82;
Memory[5481] = 8'h82;
Memory[5480] = 8'h93;
Memory[5487] = 8'h00;
Memory[5486] = 8'h62;
Memory[5485] = 8'hF2;
Memory[5484] = 8'hB3;
Memory[5491] = 8'h25;
Memory[5490] = 8'hCB;
Memory[5489] = 8'h22;
Memory[5488] = 8'h03;
Memory[5495] = 8'h00;
Memory[5494] = 8'h52;
Memory[5493] = 8'h02;
Memory[5492] = 8'h33;
Memory[5499] = 8'h00;
Memory[5498] = 8'h4B;
Memory[5497] = 8'h22;
Memory[5496] = 8'h23;
Memory[5503] = 8'h00;
Memory[5502] = 8'h0E;
Memory[5501] = 8'h8E;
Memory[5500] = 8'h13;
Memory[5507] = 8'h2C;
Memory[5506] = 8'h40;
Memory[5505] = 8'h00;
Memory[5504] = 8'h6F;
Memory[5511] = 8'h00;
Memory[5510] = 8'h82;
Memory[5509] = 8'h92;
Memory[5508] = 8'h93;
Memory[5515] = 8'h00;
Memory[5514] = 8'h92;
Memory[5513] = 8'h82;
Memory[5512] = 8'h93;
Memory[5519] = 8'h00;
Memory[5518] = 8'h62;
Memory[5517] = 8'hF2;
Memory[5516] = 8'hB3;
Memory[5523] = 8'h25;
Memory[5522] = 8'hCB;
Memory[5521] = 8'h22;
Memory[5520] = 8'h03;
Memory[5527] = 8'h00;
Memory[5526] = 8'h52;
Memory[5525] = 8'h02;
Memory[5524] = 8'h33;
Memory[5531] = 8'h00;
Memory[5530] = 8'h4B;
Memory[5529] = 8'h22;
Memory[5528] = 8'h23;
Memory[5535] = 8'h00;
Memory[5534] = 8'h0E;
Memory[5533] = 8'h8E;
Memory[5532] = 8'h13;
Memory[5539] = 8'h2C;
Memory[5538] = 8'h40;
Memory[5537] = 8'h00;
Memory[5536] = 8'h6F;
Memory[5543] = 8'h01;
Memory[5542] = 8'hF0;
Memory[5541] = 8'h01;
Memory[5540] = 8'h13;
Memory[5547] = 8'h00;
Memory[5546] = 8'h0E;
Memory[5545] = 8'h8E;
Memory[5544] = 8'h13;
Memory[5551] = 8'h0F;
Memory[5550] = 8'hF0;
Memory[5549] = 8'h01;
Memory[5548] = 8'h93;
Memory[5555] = 8'h01;
Memory[5554] = 8'h01;
Memory[5553] = 8'h91;
Memory[5552] = 8'h93;
Memory[5559] = 8'h00;
Memory[5558] = 8'h32;
Memory[5557] = 8'hF1;
Memory[5556] = 8'hB3;
Memory[5563] = 8'h01;
Memory[5562] = 8'h01;
Memory[5561] = 8'hD1;
Memory[5560] = 8'h93;
Memory[5567] = 8'h06;
Memory[5566] = 8'h40;
Memory[5565] = 8'h02;
Memory[5564] = 8'h13;
Memory[5571] = 8'h02;
Memory[5570] = 8'h41;
Memory[5569] = 8'h82;
Memory[5568] = 8'h33;
Memory[5575] = 8'h0F;
Memory[5574] = 8'hF0;
Memory[5573] = 8'h01;
Memory[5572] = 8'h93;
Memory[5579] = 8'h00;
Memory[5578] = 8'h81;
Memory[5577] = 8'h91;
Memory[5576] = 8'h93;
Memory[5583] = 8'h00;
Memory[5582] = 8'h32;
Memory[5581] = 8'hF1;
Memory[5580] = 8'hB3;
Memory[5587] = 8'h00;
Memory[5586] = 8'h81;
Memory[5585] = 8'hD1;
Memory[5584] = 8'h93;
Memory[5591] = 8'h00;
Memory[5590] = 8'hA0;
Memory[5589] = 8'h03;
Memory[5588] = 8'h13;
Memory[5595] = 8'h02;
Memory[5594] = 8'h61;
Memory[5593] = 8'h81;
Memory[5592] = 8'hB3;
Memory[5599] = 8'h00;
Memory[5598] = 8'h41;
Memory[5597] = 8'h82;
Memory[5596] = 8'h33;
Memory[5603] = 8'h0F;
Memory[5602] = 8'hF0;
Memory[5601] = 8'h01;
Memory[5600] = 8'h93;
Memory[5607] = 8'h00;
Memory[5606] = 8'h32;
Memory[5605] = 8'hF1;
Memory[5604] = 8'hB3;
Memory[5611] = 8'h00;
Memory[5610] = 8'h41;
Memory[5609] = 8'h81;
Memory[5608] = 8'hB3;
Memory[5615] = 8'h00;
Memory[5614] = 8'h3B;
Memory[5613] = 8'h2C;
Memory[5612] = 8'h23;
Memory[5619] = 8'h32;
Memory[5618] = 8'h40;
Memory[5617] = 8'h10;
Memory[5616] = 8'h6F;
Memory[5623] = 8'h01;
Memory[5622] = 8'hF0;
Memory[5621] = 8'h01;
Memory[5620] = 8'h13;
Memory[5627] = 8'h00;
Memory[5626] = 8'h0E;
Memory[5625] = 8'h8E;
Memory[5624] = 8'h13;
Memory[5631] = 8'h32;
Memory[5630] = 8'h40;
Memory[5629] = 8'h10;
Memory[5628] = 8'h6F;
Memory[5635] = 8'h02;
Memory[5634] = 8'h10;
Memory[5633] = 8'h01;
Memory[5632] = 8'h13;
Memory[5639] = 8'h18;
Memory[5638] = 8'h0B;
Memory[5637] = 8'h21;
Memory[5636] = 8'h83;
Memory[5643] = 8'h18;
Memory[5642] = 8'h4B;
Memory[5641] = 8'h22;
Memory[5640] = 8'h03;
Memory[5647] = 8'h01;
Memory[5646] = 8'hB0;
Memory[5645] = 8'h02;
Memory[5644] = 8'h93;
Memory[5651] = 8'h00;
Memory[5650] = 8'h3B;
Memory[5649] = 8'h20;
Memory[5648] = 8'h23;
Memory[5655] = 8'h00;
Memory[5654] = 8'h4B;
Memory[5653] = 8'h22;
Memory[5652] = 8'h23;
Memory[5659] = 8'h00;
Memory[5658] = 8'h5B;
Memory[5657] = 8'h24;
Memory[5656] = 8'h23;
Memory[5663] = 8'h01;
Memory[5662] = 8'hDE;
Memory[5661] = 8'h14;
Memory[5660] = 8'h63;
Memory[5667] = 8'h09;
Memory[5666] = 8'hC0;
Memory[5665] = 8'h00;
Memory[5664] = 8'h6F;
Memory[5671] = 8'h01;
Memory[5670] = 8'hDE;
Memory[5669] = 8'h42;
Memory[5668] = 8'h33;
Memory[5675] = 8'h01;
Memory[5674] = 8'h82;
Memory[5673] = 8'h71;
Memory[5672] = 8'hB3;
Memory[5679] = 8'h01;
Memory[5678] = 8'hD1;
Memory[5677] = 8'hF1;
Memory[5676] = 8'hB3;
Memory[5683] = 8'h00;
Memory[5682] = 8'h01;
Memory[5681] = 8'h84;
Memory[5680] = 8'h63;
Memory[5687] = 8'h0D;
Memory[5686] = 8'h00;
Memory[5685] = 8'h20;
Memory[5684] = 8'h6F;
Memory[5691] = 8'hFF;
Memory[5690] = 8'hF2;
Memory[5689] = 8'h71;
Memory[5688] = 8'h93;
Memory[5695] = 8'h01;
Memory[5694] = 8'hD1;
Memory[5693] = 8'hF1;
Memory[5692] = 8'hB3;
Memory[5699] = 8'h00;
Memory[5698] = 8'h01;
Memory[5697] = 8'h94;
Memory[5696] = 8'h63;
Memory[5703] = 8'h2C;
Memory[5702] = 8'h40;
Memory[5701] = 8'h00;
Memory[5700] = 8'h6F;
Memory[5707] = 8'h10;
Memory[5706] = 8'h01;
Memory[5705] = 8'hF2;
Memory[5704] = 8'h13;
Memory[5711] = 8'h00;
Memory[5710] = 8'h02;
Memory[5709] = 8'h18;
Memory[5708] = 8'h63;
Memory[5715] = 8'h00;
Memory[5714] = 8'h41;
Memory[5713] = 8'hF2;
Memory[5712] = 8'h13;
Memory[5719] = 8'h00;
Memory[5718] = 8'h02;
Memory[5717] = 8'h1A;
Memory[5716] = 8'h63;
Memory[5723] = 8'h2C;
Memory[5722] = 8'h40;
Memory[5721] = 8'h00;
Memory[5720] = 8'h6F;
Memory[5727] = 8'h01;
Memory[5726] = 8'h30;
Memory[5725] = 8'h01;
Memory[5724] = 8'h13;
Memory[5731] = 8'h00;
Memory[5730] = 8'h0E;
Memory[5729] = 8'h8E;
Memory[5728] = 8'h13;
Memory[5735] = 8'h37;
Memory[5734] = 8'h50;
Memory[5733] = 8'h00;
Memory[5732] = 8'h6F;
Memory[5739] = 8'h01;
Memory[5738] = 8'hF0;
Memory[5737] = 8'h01;
Memory[5736] = 8'h13;
Memory[5743] = 8'h00;
Memory[5742] = 8'h0E;
Memory[5741] = 8'h8E;
Memory[5740] = 8'h13;
Memory[5747] = 8'h32;
Memory[5746] = 8'h40;
Memory[5745] = 8'h10;
Memory[5744] = 8'h6F;
Memory[5751] = 8'h02;
Memory[5750] = 8'h50;
Memory[5749] = 8'h01;
Memory[5748] = 8'h13;
Memory[5755] = 8'h1C;
Memory[5754] = 8'h8B;
Memory[5753] = 8'h21;
Memory[5752] = 8'h83;
Memory[5759] = 8'h1C;
Memory[5758] = 8'hCB;
Memory[5757] = 8'h22;
Memory[5756] = 8'h03;
Memory[5763] = 8'h00;
Memory[5762] = 8'hC0;
Memory[5761] = 8'h02;
Memory[5760] = 8'h93;
Memory[5767] = 8'h00;
Memory[5766] = 8'h3B;
Memory[5765] = 8'h20;
Memory[5764] = 8'h23;
Memory[5771] = 8'h00;
Memory[5770] = 8'h4B;
Memory[5769] = 8'h22;
Memory[5768] = 8'h23;
Memory[5775] = 8'h00;
Memory[5774] = 8'h5B;
Memory[5773] = 8'h24;
Memory[5772] = 8'h23;
Memory[5779] = 8'h01;
Memory[5778] = 8'hDE;
Memory[5777] = 8'h14;
Memory[5776] = 8'h63;
Memory[5783] = 8'h09;
Memory[5782] = 8'hC0;
Memory[5781] = 8'h00;
Memory[5780] = 8'h6F;
Memory[5787] = 8'h01;
Memory[5786] = 8'hDE;
Memory[5785] = 8'h42;
Memory[5784] = 8'h33;
Memory[5791] = 8'h01;
Memory[5790] = 8'h82;
Memory[5789] = 8'h71;
Memory[5788] = 8'hB3;
Memory[5795] = 8'h01;
Memory[5794] = 8'hD1;
Memory[5793] = 8'hF1;
Memory[5792] = 8'hB3;
Memory[5799] = 8'h00;
Memory[5798] = 8'h01;
Memory[5797] = 8'h84;
Memory[5796] = 8'h63;
Memory[5803] = 8'h0D;
Memory[5802] = 8'h00;
Memory[5801] = 8'h20;
Memory[5800] = 8'h6F;
Memory[5807] = 8'hFF;
Memory[5806] = 8'hF2;
Memory[5805] = 8'h71;
Memory[5804] = 8'h93;
Memory[5811] = 8'h01;
Memory[5810] = 8'hD1;
Memory[5809] = 8'hF1;
Memory[5808] = 8'hB3;
Memory[5815] = 8'h00;
Memory[5814] = 8'h01;
Memory[5813] = 8'h94;
Memory[5812] = 8'h63;
Memory[5819] = 8'h2C;
Memory[5818] = 8'h40;
Memory[5817] = 8'h00;
Memory[5816] = 8'h6F;
Memory[5823] = 8'h04;
Memory[5822] = 8'h01;
Memory[5821] = 8'hF2;
Memory[5820] = 8'h13;
Memory[5827] = 8'h00;
Memory[5826] = 8'h02;
Memory[5825] = 8'h1C;
Memory[5824] = 8'h63;
Memory[5831] = 8'h00;
Memory[5830] = 8'h41;
Memory[5829] = 8'hF2;
Memory[5828] = 8'h13;
Memory[5835] = 8'h00;
Memory[5834] = 8'h02;
Memory[5833] = 8'h1E;
Memory[5832] = 8'h63;
Memory[5839] = 8'h00;
Memory[5838] = 8'h11;
Memory[5837] = 8'hF2;
Memory[5836] = 8'h13;
Memory[5843] = 8'h02;
Memory[5842] = 8'h02;
Memory[5841] = 8'h10;
Memory[5840] = 8'h63;
Memory[5847] = 8'h2C;
Memory[5846] = 8'h40;
Memory[5845] = 8'h00;
Memory[5844] = 8'h6F;
Memory[5851] = 8'h02;
Memory[5850] = 8'h60;
Memory[5849] = 8'h01;
Memory[5848] = 8'h13;
Memory[5855] = 8'h00;
Memory[5854] = 8'h0E;
Memory[5853] = 8'h8E;
Memory[5852] = 8'h13;
Memory[5859] = 8'h6F;
Memory[5858] = 8'hC0;
Memory[5857] = 8'h10;
Memory[5856] = 8'h6F;
Memory[5863] = 8'h02;
Memory[5862] = 8'h90;
Memory[5861] = 8'h01;
Memory[5860] = 8'h13;
Memory[5867] = 8'h00;
Memory[5866] = 8'h0E;
Memory[5865] = 8'h8E;
Memory[5864] = 8'h13;
Memory[5871] = 8'h0B;
Memory[5870] = 8'h50;
Memory[5869] = 8'h10;
Memory[5868] = 8'h6F;
Memory[5875] = 8'h00;
Memory[5874] = 8'h80;
Memory[5873] = 8'h01;
Memory[5872] = 8'h13;
Memory[5879] = 8'h00;
Memory[5878] = 8'h0E;
Memory[5877] = 8'h8E;
Memory[5876] = 8'h13;
Memory[5883] = 8'h6A;
Memory[5882] = 8'h80;
Memory[5881] = 8'h00;
Memory[5880] = 8'h6F;
Memory[5887] = 8'h02;
Memory[5886] = 8'h60;
Memory[5885] = 8'h01;
Memory[5884] = 8'h13;
Memory[5891] = 8'h1D;
Memory[5890] = 8'h0B;
Memory[5889] = 8'h21;
Memory[5888] = 8'h83;
Memory[5895] = 8'h1D;
Memory[5894] = 8'h4B;
Memory[5893] = 8'h22;
Memory[5892] = 8'h03;
Memory[5899] = 8'h00;
Memory[5898] = 8'hB0;
Memory[5897] = 8'h02;
Memory[5896] = 8'h93;
Memory[5903] = 8'h00;
Memory[5902] = 8'h3B;
Memory[5901] = 8'h20;
Memory[5900] = 8'h23;
Memory[5907] = 8'h00;
Memory[5906] = 8'h4B;
Memory[5905] = 8'h22;
Memory[5904] = 8'h23;
Memory[5911] = 8'h00;
Memory[5910] = 8'h5B;
Memory[5909] = 8'h24;
Memory[5908] = 8'h23;
Memory[5915] = 8'h01;
Memory[5914] = 8'hDE;
Memory[5913] = 8'h14;
Memory[5912] = 8'h63;
Memory[5919] = 8'h09;
Memory[5918] = 8'hC0;
Memory[5917] = 8'h00;
Memory[5916] = 8'h6F;
Memory[5923] = 8'h01;
Memory[5922] = 8'hDE;
Memory[5921] = 8'h42;
Memory[5920] = 8'h33;
Memory[5927] = 8'h01;
Memory[5926] = 8'h82;
Memory[5925] = 8'h71;
Memory[5924] = 8'hB3;
Memory[5931] = 8'h01;
Memory[5930] = 8'hD1;
Memory[5929] = 8'hF1;
Memory[5928] = 8'hB3;
Memory[5935] = 8'h00;
Memory[5934] = 8'h01;
Memory[5933] = 8'h84;
Memory[5932] = 8'h63;
Memory[5939] = 8'h0D;
Memory[5938] = 8'h00;
Memory[5937] = 8'h20;
Memory[5936] = 8'h6F;
Memory[5943] = 8'hFF;
Memory[5942] = 8'hF2;
Memory[5941] = 8'h71;
Memory[5940] = 8'h93;
Memory[5947] = 8'h01;
Memory[5946] = 8'hD1;
Memory[5945] = 8'hF1;
Memory[5944] = 8'hB3;
Memory[5951] = 8'h00;
Memory[5950] = 8'h01;
Memory[5949] = 8'h94;
Memory[5948] = 8'h63;
Memory[5955] = 8'h2C;
Memory[5954] = 8'h40;
Memory[5953] = 8'h00;
Memory[5952] = 8'h6F;
Memory[5959] = 8'h10;
Memory[5958] = 8'h01;
Memory[5957] = 8'hF2;
Memory[5956] = 8'h13;
Memory[5963] = 8'h00;
Memory[5962] = 8'h02;
Memory[5961] = 8'h1C;
Memory[5960] = 8'h63;
Memory[5967] = 8'h00;
Memory[5966] = 8'h41;
Memory[5965] = 8'hF2;
Memory[5964] = 8'h13;
Memory[5971] = 8'h00;
Memory[5970] = 8'h02;
Memory[5969] = 8'h1E;
Memory[5968] = 8'h63;
Memory[5975] = 8'h00;
Memory[5974] = 8'h11;
Memory[5973] = 8'hF2;
Memory[5972] = 8'h13;
Memory[5979] = 8'h02;
Memory[5978] = 8'h02;
Memory[5977] = 8'h10;
Memory[5976] = 8'h63;
Memory[5983] = 8'h2C;
Memory[5982] = 8'h40;
Memory[5981] = 8'h00;
Memory[5980] = 8'h6F;
Memory[5987] = 8'h02;
Memory[5986] = 8'h50;
Memory[5985] = 8'h01;
Memory[5984] = 8'h13;
Memory[5991] = 8'h00;
Memory[5990] = 8'h0E;
Memory[5989] = 8'h8E;
Memory[5988] = 8'h13;
Memory[5995] = 8'h67;
Memory[5994] = 8'h40;
Memory[5993] = 8'h10;
Memory[5992] = 8'h6F;
Memory[5999] = 8'h02;
Memory[5998] = 8'h70;
Memory[5997] = 8'h01;
Memory[5996] = 8'h13;
Memory[6003] = 8'h00;
Memory[6002] = 8'h0E;
Memory[6001] = 8'h8E;
Memory[6000] = 8'h13;
Memory[6007] = 8'h78;
Memory[6006] = 8'h40;
Memory[6005] = 8'h10;
Memory[6004] = 8'h6F;
Memory[6011] = 8'h00;
Memory[6010] = 8'h80;
Memory[6009] = 8'h01;
Memory[6008] = 8'h13;
Memory[6015] = 8'h00;
Memory[6014] = 8'h0E;
Memory[6013] = 8'h8E;
Memory[6012] = 8'h13;
Memory[6019] = 8'h6A;
Memory[6018] = 8'h80;
Memory[6017] = 8'h00;
Memory[6016] = 8'h6F;
Memory[6023] = 8'h02;
Memory[6022] = 8'h70;
Memory[6021] = 8'h01;
Memory[6020] = 8'h13;
Memory[6027] = 8'h1D;
Memory[6026] = 8'h8B;
Memory[6025] = 8'h21;
Memory[6024] = 8'h83;
Memory[6031] = 8'h1D;
Memory[6030] = 8'hCB;
Memory[6029] = 8'h22;
Memory[6028] = 8'h03;
Memory[6035] = 8'h00;
Memory[6034] = 8'hE0;
Memory[6033] = 8'h02;
Memory[6032] = 8'h93;
Memory[6039] = 8'h00;
Memory[6038] = 8'h3B;
Memory[6037] = 8'h20;
Memory[6036] = 8'h23;
Memory[6043] = 8'h00;
Memory[6042] = 8'h4B;
Memory[6041] = 8'h22;
Memory[6040] = 8'h23;
Memory[6047] = 8'h00;
Memory[6046] = 8'h5B;
Memory[6045] = 8'h24;
Memory[6044] = 8'h23;
Memory[6051] = 8'h01;
Memory[6050] = 8'hDE;
Memory[6049] = 8'h14;
Memory[6048] = 8'h63;
Memory[6055] = 8'h09;
Memory[6054] = 8'hC0;
Memory[6053] = 8'h00;
Memory[6052] = 8'h6F;
Memory[6059] = 8'h01;
Memory[6058] = 8'hDE;
Memory[6057] = 8'h42;
Memory[6056] = 8'h33;
Memory[6063] = 8'h01;
Memory[6062] = 8'h82;
Memory[6061] = 8'h71;
Memory[6060] = 8'hB3;
Memory[6067] = 8'h01;
Memory[6066] = 8'hD1;
Memory[6065] = 8'hF1;
Memory[6064] = 8'hB3;
Memory[6071] = 8'h00;
Memory[6070] = 8'h01;
Memory[6069] = 8'h84;
Memory[6068] = 8'h63;
Memory[6075] = 8'h0D;
Memory[6074] = 8'h00;
Memory[6073] = 8'h20;
Memory[6072] = 8'h6F;
Memory[6079] = 8'hFF;
Memory[6078] = 8'hF2;
Memory[6077] = 8'h71;
Memory[6076] = 8'h93;
Memory[6083] = 8'h01;
Memory[6082] = 8'hD1;
Memory[6081] = 8'hF1;
Memory[6080] = 8'hB3;
Memory[6087] = 8'h00;
Memory[6086] = 8'h01;
Memory[6085] = 8'h94;
Memory[6084] = 8'h63;
Memory[6091] = 8'h2C;
Memory[6090] = 8'h40;
Memory[6089] = 8'h00;
Memory[6088] = 8'h6F;
Memory[6095] = 8'h01;
Memory[6094] = 8'h01;
Memory[6093] = 8'hF2;
Memory[6092] = 8'h13;
Memory[6099] = 8'h00;
Memory[6098] = 8'h02;
Memory[6097] = 8'h1C;
Memory[6096] = 8'h63;
Memory[6103] = 8'h00;
Memory[6102] = 8'h41;
Memory[6101] = 8'hF2;
Memory[6100] = 8'h13;
Memory[6107] = 8'h00;
Memory[6106] = 8'h02;
Memory[6105] = 8'h1E;
Memory[6104] = 8'h63;
Memory[6111] = 8'h00;
Memory[6110] = 8'h11;
Memory[6109] = 8'hF2;
Memory[6108] = 8'h13;
Memory[6115] = 8'h02;
Memory[6114] = 8'h02;
Memory[6113] = 8'h18;
Memory[6112] = 8'h63;
Memory[6119] = 8'h2C;
Memory[6118] = 8'h40;
Memory[6117] = 8'h00;
Memory[6116] = 8'h6F;
Memory[6123] = 8'h02;
Memory[6122] = 8'h80;
Memory[6121] = 8'h01;
Memory[6120] = 8'h13;
Memory[6127] = 8'h00;
Memory[6126] = 8'h0E;
Memory[6125] = 8'h8E;
Memory[6124] = 8'h13;
Memory[6131] = 8'h01;
Memory[6130] = 8'hD0;
Memory[6129] = 8'h10;
Memory[6128] = 8'h6F;
Memory[6135] = 8'h02;
Memory[6134] = 8'hB0;
Memory[6133] = 8'h01;
Memory[6132] = 8'h13;
Memory[6139] = 8'h00;
Memory[6138] = 8'h0E;
Memory[6137] = 8'h8E;
Memory[6136] = 8'h13;
Memory[6143] = 8'h00;
Memory[6142] = 8'h30;
Memory[6141] = 8'h01;
Memory[6140] = 8'h93;
Memory[6147] = 8'h26;
Memory[6146] = 8'h3B;
Memory[6145] = 8'h20;
Memory[6144] = 8'h23;
Memory[6151] = 8'h08;
Memory[6150] = 8'h0B;
Memory[6149] = 8'h2E;
Memory[6148] = 8'h23;
Memory[6155] = 8'h05;
Memory[6154] = 8'hFB;
Memory[6153] = 8'h28;
Memory[6152] = 8'h23;
Memory[6159] = 8'h1E;
Memory[6158] = 8'h50;
Memory[6157] = 8'h10;
Memory[6156] = 8'h6F;
Memory[6163] = 8'h02;
Memory[6162] = 8'h60;
Memory[6161] = 8'h01;
Memory[6160] = 8'h13;
Memory[6167] = 8'h00;
Memory[6166] = 8'h0E;
Memory[6165] = 8'h8E;
Memory[6164] = 8'h13;
Memory[6171] = 8'h6F;
Memory[6170] = 8'hC0;
Memory[6169] = 8'h10;
Memory[6168] = 8'h6F;
Memory[6175] = 8'h02;
Memory[6174] = 8'h80;
Memory[6173] = 8'h01;
Memory[6172] = 8'h13;
Memory[6179] = 8'h1E;
Memory[6178] = 8'h0B;
Memory[6177] = 8'h21;
Memory[6176] = 8'h83;
Memory[6183] = 8'h1E;
Memory[6182] = 8'h4B;
Memory[6181] = 8'h22;
Memory[6180] = 8'h03;
Memory[6187] = 8'h01;
Memory[6186] = 8'h10;
Memory[6185] = 8'h02;
Memory[6184] = 8'h93;
Memory[6191] = 8'h00;
Memory[6190] = 8'h3B;
Memory[6189] = 8'h20;
Memory[6188] = 8'h23;
Memory[6195] = 8'h00;
Memory[6194] = 8'h4B;
Memory[6193] = 8'h22;
Memory[6192] = 8'h23;
Memory[6199] = 8'h00;
Memory[6198] = 8'h5B;
Memory[6197] = 8'h24;
Memory[6196] = 8'h23;
Memory[6203] = 8'h01;
Memory[6202] = 8'hDE;
Memory[6201] = 8'h14;
Memory[6200] = 8'h63;
Memory[6207] = 8'h09;
Memory[6206] = 8'hC0;
Memory[6205] = 8'h00;
Memory[6204] = 8'h6F;
Memory[6211] = 8'h01;
Memory[6210] = 8'hDE;
Memory[6209] = 8'h42;
Memory[6208] = 8'h33;
Memory[6215] = 8'h01;
Memory[6214] = 8'h82;
Memory[6213] = 8'h71;
Memory[6212] = 8'hB3;
Memory[6219] = 8'h01;
Memory[6218] = 8'hD1;
Memory[6217] = 8'hF1;
Memory[6216] = 8'hB3;
Memory[6223] = 8'h00;
Memory[6222] = 8'h01;
Memory[6221] = 8'h84;
Memory[6220] = 8'h63;
Memory[6227] = 8'h0D;
Memory[6226] = 8'h00;
Memory[6225] = 8'h20;
Memory[6224] = 8'h6F;
Memory[6231] = 8'hFF;
Memory[6230] = 8'hF2;
Memory[6229] = 8'h71;
Memory[6228] = 8'h93;
Memory[6235] = 8'h01;
Memory[6234] = 8'hD1;
Memory[6233] = 8'hF1;
Memory[6232] = 8'hB3;
Memory[6239] = 8'h00;
Memory[6238] = 8'h01;
Memory[6237] = 8'h94;
Memory[6236] = 8'h63;
Memory[6243] = 8'h2C;
Memory[6242] = 8'h40;
Memory[6241] = 8'h00;
Memory[6240] = 8'h6F;
Memory[6247] = 8'h40;
Memory[6246] = 8'h01;
Memory[6245] = 8'hF2;
Memory[6244] = 8'h13;
Memory[6251] = 8'h00;
Memory[6250] = 8'h02;
Memory[6249] = 8'h1C;
Memory[6248] = 8'h63;
Memory[6255] = 8'h00;
Memory[6254] = 8'h41;
Memory[6253] = 8'hF2;
Memory[6252] = 8'h13;
Memory[6259] = 8'h00;
Memory[6258] = 8'h02;
Memory[6257] = 8'h1E;
Memory[6256] = 8'h63;
Memory[6263] = 8'h00;
Memory[6262] = 8'h11;
Memory[6261] = 8'hF2;
Memory[6260] = 8'h13;
Memory[6267] = 8'h02;
Memory[6266] = 8'h02;
Memory[6265] = 8'h18;
Memory[6264] = 8'h63;
Memory[6271] = 8'h2C;
Memory[6270] = 8'h40;
Memory[6269] = 8'h00;
Memory[6268] = 8'h6F;
Memory[6275] = 8'h02;
Memory[6274] = 8'h70;
Memory[6273] = 8'h01;
Memory[6272] = 8'h13;
Memory[6279] = 8'h00;
Memory[6278] = 8'h0E;
Memory[6277] = 8'h8E;
Memory[6276] = 8'h13;
Memory[6283] = 8'h78;
Memory[6282] = 8'h40;
Memory[6281] = 8'h10;
Memory[6280] = 8'h6F;
Memory[6287] = 8'h02;
Memory[6286] = 8'hB0;
Memory[6285] = 8'h01;
Memory[6284] = 8'h13;
Memory[6291] = 8'h00;
Memory[6290] = 8'h0E;
Memory[6289] = 8'h8E;
Memory[6288] = 8'h13;
Memory[6295] = 8'h00;
Memory[6294] = 8'h40;
Memory[6293] = 8'h01;
Memory[6292] = 8'h93;
Memory[6299] = 8'h26;
Memory[6298] = 8'h3B;
Memory[6297] = 8'h20;
Memory[6296] = 8'h23;
Memory[6303] = 8'h08;
Memory[6302] = 8'h0B;
Memory[6301] = 8'h2E;
Memory[6300] = 8'h23;
Memory[6307] = 8'h05;
Memory[6306] = 8'hFB;
Memory[6305] = 8'h28;
Memory[6304] = 8'h23;
Memory[6311] = 8'h1E;
Memory[6310] = 8'h50;
Memory[6309] = 8'h10;
Memory[6308] = 8'h6F;
Memory[6315] = 8'h02;
Memory[6314] = 8'h60;
Memory[6313] = 8'h01;
Memory[6312] = 8'h13;
Memory[6319] = 8'h00;
Memory[6318] = 8'h0E;
Memory[6317] = 8'h8E;
Memory[6316] = 8'h13;
Memory[6323] = 8'h6F;
Memory[6322] = 8'hC0;
Memory[6321] = 8'h10;
Memory[6320] = 8'h6F;
Memory[6327] = 8'h02;
Memory[6326] = 8'h90;
Memory[6325] = 8'h01;
Memory[6324] = 8'h13;
Memory[6331] = 8'h1D;
Memory[6330] = 8'h8B;
Memory[6329] = 8'h21;
Memory[6328] = 8'h83;
Memory[6335] = 8'h1D;
Memory[6334] = 8'hCB;
Memory[6333] = 8'h22;
Memory[6332] = 8'h03;
Memory[6339] = 8'h00;
Memory[6338] = 8'hE0;
Memory[6337] = 8'h02;
Memory[6336] = 8'h93;
Memory[6343] = 8'h00;
Memory[6342] = 8'h3B;
Memory[6341] = 8'h20;
Memory[6340] = 8'h23;
Memory[6347] = 8'h00;
Memory[6346] = 8'h4B;
Memory[6345] = 8'h22;
Memory[6344] = 8'h23;
Memory[6351] = 8'h00;
Memory[6350] = 8'h5B;
Memory[6349] = 8'h24;
Memory[6348] = 8'h23;
Memory[6355] = 8'h01;
Memory[6354] = 8'hDE;
Memory[6353] = 8'h14;
Memory[6352] = 8'h63;
Memory[6359] = 8'h09;
Memory[6358] = 8'hC0;
Memory[6357] = 8'h00;
Memory[6356] = 8'h6F;
Memory[6363] = 8'h01;
Memory[6362] = 8'hDE;
Memory[6361] = 8'h42;
Memory[6360] = 8'h33;
Memory[6367] = 8'h01;
Memory[6366] = 8'h82;
Memory[6365] = 8'h71;
Memory[6364] = 8'hB3;
Memory[6371] = 8'h01;
Memory[6370] = 8'hD1;
Memory[6369] = 8'hF1;
Memory[6368] = 8'hB3;
Memory[6375] = 8'h00;
Memory[6374] = 8'h01;
Memory[6373] = 8'h84;
Memory[6372] = 8'h63;
Memory[6379] = 8'h0D;
Memory[6378] = 8'h00;
Memory[6377] = 8'h20;
Memory[6376] = 8'h6F;
Memory[6383] = 8'hFF;
Memory[6382] = 8'hF2;
Memory[6381] = 8'h71;
Memory[6380] = 8'h93;
Memory[6387] = 8'h01;
Memory[6386] = 8'hD1;
Memory[6385] = 8'hF1;
Memory[6384] = 8'hB3;
Memory[6391] = 8'h00;
Memory[6390] = 8'h01;
Memory[6389] = 8'h94;
Memory[6388] = 8'h63;
Memory[6395] = 8'h2C;
Memory[6394] = 8'h40;
Memory[6393] = 8'h00;
Memory[6392] = 8'h6F;
Memory[6399] = 8'h01;
Memory[6398] = 8'h01;
Memory[6397] = 8'hF2;
Memory[6396] = 8'h13;
Memory[6403] = 8'h00;
Memory[6402] = 8'h02;
Memory[6401] = 8'h1C;
Memory[6400] = 8'h63;
Memory[6407] = 8'h00;
Memory[6406] = 8'h41;
Memory[6405] = 8'hF2;
Memory[6404] = 8'h13;
Memory[6411] = 8'h00;
Memory[6410] = 8'h02;
Memory[6409] = 8'h1E;
Memory[6408] = 8'h63;
Memory[6415] = 8'h00;
Memory[6414] = 8'h11;
Memory[6413] = 8'hF2;
Memory[6412] = 8'h13;
Memory[6419] = 8'h02;
Memory[6418] = 8'h02;
Memory[6417] = 8'h18;
Memory[6416] = 8'h63;
Memory[6423] = 8'h2C;
Memory[6422] = 8'h40;
Memory[6421] = 8'h00;
Memory[6420] = 8'h6F;
Memory[6427] = 8'h02;
Memory[6426] = 8'hA0;
Memory[6425] = 8'h01;
Memory[6424] = 8'h13;
Memory[6431] = 8'h00;
Memory[6430] = 8'h0E;
Memory[6429] = 8'h8E;
Memory[6428] = 8'h13;
Memory[6435] = 8'h14;
Memory[6434] = 8'hD0;
Memory[6433] = 8'h10;
Memory[6432] = 8'h6F;
Memory[6439] = 8'h02;
Memory[6438] = 8'hB0;
Memory[6437] = 8'h01;
Memory[6436] = 8'h13;
Memory[6443] = 8'h00;
Memory[6442] = 8'h0E;
Memory[6441] = 8'h8E;
Memory[6440] = 8'h13;
Memory[6447] = 8'h00;
Memory[6446] = 8'h10;
Memory[6445] = 8'h01;
Memory[6444] = 8'h93;
Memory[6451] = 8'h26;
Memory[6450] = 8'h3B;
Memory[6449] = 8'h20;
Memory[6448] = 8'h23;
Memory[6455] = 8'h08;
Memory[6454] = 8'h0B;
Memory[6453] = 8'h2E;
Memory[6452] = 8'h23;
Memory[6459] = 8'h05;
Memory[6458] = 8'hFB;
Memory[6457] = 8'h28;
Memory[6456] = 8'h23;
Memory[6463] = 8'h1E;
Memory[6462] = 8'h50;
Memory[6461] = 8'h10;
Memory[6460] = 8'h6F;
Memory[6467] = 8'h02;
Memory[6466] = 8'h50;
Memory[6465] = 8'h01;
Memory[6464] = 8'h13;
Memory[6471] = 8'h00;
Memory[6470] = 8'h0E;
Memory[6469] = 8'h8E;
Memory[6468] = 8'h13;
Memory[6475] = 8'h67;
Memory[6474] = 8'h40;
Memory[6473] = 8'h10;
Memory[6472] = 8'h6F;
Memory[6479] = 8'h02;
Memory[6478] = 8'hA0;
Memory[6477] = 8'h01;
Memory[6476] = 8'h13;
Memory[6483] = 8'h1E;
Memory[6482] = 8'h0B;
Memory[6481] = 8'h21;
Memory[6480] = 8'h83;
Memory[6487] = 8'h1E;
Memory[6486] = 8'h4B;
Memory[6485] = 8'h22;
Memory[6484] = 8'h03;
Memory[6491] = 8'h01;
Memory[6490] = 8'h10;
Memory[6489] = 8'h02;
Memory[6488] = 8'h93;
Memory[6495] = 8'h00;
Memory[6494] = 8'h3B;
Memory[6493] = 8'h20;
Memory[6492] = 8'h23;
Memory[6499] = 8'h00;
Memory[6498] = 8'h4B;
Memory[6497] = 8'h22;
Memory[6496] = 8'h23;
Memory[6503] = 8'h00;
Memory[6502] = 8'h5B;
Memory[6501] = 8'h24;
Memory[6500] = 8'h23;
Memory[6507] = 8'h01;
Memory[6506] = 8'hDE;
Memory[6505] = 8'h14;
Memory[6504] = 8'h63;
Memory[6511] = 8'h09;
Memory[6510] = 8'hC0;
Memory[6509] = 8'h00;
Memory[6508] = 8'h6F;
Memory[6515] = 8'h01;
Memory[6514] = 8'hDE;
Memory[6513] = 8'h42;
Memory[6512] = 8'h33;
Memory[6519] = 8'h01;
Memory[6518] = 8'h82;
Memory[6517] = 8'h71;
Memory[6516] = 8'hB3;
Memory[6523] = 8'h01;
Memory[6522] = 8'hD1;
Memory[6521] = 8'hF1;
Memory[6520] = 8'hB3;
Memory[6527] = 8'h00;
Memory[6526] = 8'h01;
Memory[6525] = 8'h84;
Memory[6524] = 8'h63;
Memory[6531] = 8'h0D;
Memory[6530] = 8'h00;
Memory[6529] = 8'h20;
Memory[6528] = 8'h6F;
Memory[6535] = 8'hFF;
Memory[6534] = 8'hF2;
Memory[6533] = 8'h71;
Memory[6532] = 8'h93;
Memory[6539] = 8'h01;
Memory[6538] = 8'hD1;
Memory[6537] = 8'hF1;
Memory[6536] = 8'hB3;
Memory[6543] = 8'h00;
Memory[6542] = 8'h01;
Memory[6541] = 8'h94;
Memory[6540] = 8'h63;
Memory[6547] = 8'h2C;
Memory[6546] = 8'h40;
Memory[6545] = 8'h00;
Memory[6544] = 8'h6F;
Memory[6551] = 8'h40;
Memory[6550] = 8'h01;
Memory[6549] = 8'hF2;
Memory[6548] = 8'h13;
Memory[6555] = 8'h00;
Memory[6554] = 8'h02;
Memory[6553] = 8'h1C;
Memory[6552] = 8'h63;
Memory[6559] = 8'h00;
Memory[6558] = 8'h41;
Memory[6557] = 8'hF2;
Memory[6556] = 8'h13;
Memory[6563] = 8'h00;
Memory[6562] = 8'h02;
Memory[6561] = 8'h1E;
Memory[6560] = 8'h63;
Memory[6567] = 8'h00;
Memory[6566] = 8'h11;
Memory[6565] = 8'hF2;
Memory[6564] = 8'h13;
Memory[6571] = 8'h02;
Memory[6570] = 8'h02;
Memory[6569] = 8'h18;
Memory[6568] = 8'h63;
Memory[6575] = 8'h2C;
Memory[6574] = 8'h40;
Memory[6573] = 8'h00;
Memory[6572] = 8'h6F;
Memory[6579] = 8'h02;
Memory[6578] = 8'h90;
Memory[6577] = 8'h01;
Memory[6576] = 8'h13;
Memory[6583] = 8'h00;
Memory[6582] = 8'h0E;
Memory[6581] = 8'h8E;
Memory[6580] = 8'h13;
Memory[6587] = 8'h0B;
Memory[6586] = 8'h50;
Memory[6585] = 8'h10;
Memory[6584] = 8'h6F;
Memory[6591] = 8'h02;
Memory[6590] = 8'hB0;
Memory[6589] = 8'h01;
Memory[6588] = 8'h13;
Memory[6595] = 8'h00;
Memory[6594] = 8'h0E;
Memory[6593] = 8'h8E;
Memory[6592] = 8'h13;
Memory[6599] = 8'h00;
Memory[6598] = 8'h20;
Memory[6597] = 8'h01;
Memory[6596] = 8'h93;
Memory[6603] = 8'h26;
Memory[6602] = 8'h3B;
Memory[6601] = 8'h20;
Memory[6600] = 8'h23;
Memory[6607] = 8'h08;
Memory[6606] = 8'h0B;
Memory[6605] = 8'h2E;
Memory[6604] = 8'h23;
Memory[6611] = 8'h05;
Memory[6610] = 8'hFB;
Memory[6609] = 8'h28;
Memory[6608] = 8'h23;
Memory[6615] = 8'h1E;
Memory[6614] = 8'h50;
Memory[6613] = 8'h10;
Memory[6612] = 8'h6F;
Memory[6619] = 8'h02;
Memory[6618] = 8'h50;
Memory[6617] = 8'h01;
Memory[6616] = 8'h13;
Memory[6623] = 8'h00;
Memory[6622] = 8'h0E;
Memory[6621] = 8'h8E;
Memory[6620] = 8'h13;
Memory[6627] = 8'h67;
Memory[6626] = 8'h40;
Memory[6625] = 8'h10;
Memory[6624] = 8'h6F;
Memory[6631] = 8'h02;
Memory[6630] = 8'hB0;
Memory[6629] = 8'h01;
Memory[6628] = 8'h13;
Memory[6635] = 8'h01;
Memory[6634] = 8'h00;
Memory[6633] = 8'h01;
Memory[6632] = 8'h93;
Memory[6639] = 8'h00;
Memory[6638] = 8'h3B;
Memory[6637] = 8'h24;
Memory[6636] = 8'h23;
Memory[6643] = 8'h01;
Memory[6642] = 8'hDE;
Memory[6641] = 8'h14;
Memory[6640] = 8'h63;
Memory[6647] = 8'h09;
Memory[6646] = 8'hC0;
Memory[6645] = 8'h00;
Memory[6644] = 8'h6F;
Memory[6651] = 8'h01;
Memory[6650] = 8'hDE;
Memory[6649] = 8'h42;
Memory[6648] = 8'h33;
Memory[6655] = 8'h01;
Memory[6654] = 8'h82;
Memory[6653] = 8'h71;
Memory[6652] = 8'hB3;
Memory[6659] = 8'h01;
Memory[6658] = 8'hD1;
Memory[6657] = 8'hF1;
Memory[6656] = 8'hB3;
Memory[6663] = 8'h00;
Memory[6662] = 8'h01;
Memory[6661] = 8'h84;
Memory[6660] = 8'h63;
Memory[6667] = 8'h0D;
Memory[6666] = 8'h00;
Memory[6665] = 8'h20;
Memory[6664] = 8'h6F;
Memory[6671] = 8'h01;
Memory[6670] = 8'h72;
Memory[6669] = 8'h71;
Memory[6668] = 8'hB3;
Memory[6675] = 8'h01;
Memory[6674] = 8'hD1;
Memory[6673] = 8'hF1;
Memory[6672] = 8'hB3;
Memory[6679] = 8'h00;
Memory[6678] = 8'h01;
Memory[6677] = 8'h8C;
Memory[6676] = 8'h63;
Memory[6683] = 8'h02;
Memory[6682] = 8'hE0;
Memory[6681] = 8'h01;
Memory[6680] = 8'h13;
Memory[6687] = 8'h00;
Memory[6686] = 8'h0E;
Memory[6685] = 8'h8E;
Memory[6684] = 8'h13;
Memory[6691] = 8'h00;
Memory[6690] = 8'h0F;
Memory[6689] = 8'h81;
Memory[6688] = 8'h93;
Memory[6695] = 8'h08;
Memory[6694] = 8'h3B;
Memory[6693] = 8'h2E;
Memory[6692] = 8'h23;
Memory[6699] = 8'h23;
Memory[6698] = 8'h10;
Memory[6697] = 8'h10;
Memory[6696] = 8'h6F;
Memory[6703] = 8'h2C;
Memory[6702] = 8'h40;
Memory[6701] = 8'h00;
Memory[6700] = 8'h6F;
Memory[6707] = 8'h02;
Memory[6706] = 8'hE0;
Memory[6705] = 8'h01;
Memory[6704] = 8'h13;
Memory[6711] = 8'h1F;
Memory[6710] = 8'h8B;
Memory[6709] = 8'h21;
Memory[6708] = 8'h83;
Memory[6715] = 8'h1F;
Memory[6714] = 8'hCB;
Memory[6713] = 8'h22;
Memory[6712] = 8'h03;
Memory[6719] = 8'h01;
Memory[6718] = 8'h80;
Memory[6717] = 8'h02;
Memory[6716] = 8'h93;
Memory[6723] = 8'h00;
Memory[6722] = 8'h3B;
Memory[6721] = 8'h20;
Memory[6720] = 8'h23;
Memory[6727] = 8'h00;
Memory[6726] = 8'h4B;
Memory[6725] = 8'h22;
Memory[6724] = 8'h23;
Memory[6731] = 8'h00;
Memory[6730] = 8'h5B;
Memory[6729] = 8'h24;
Memory[6728] = 8'h23;
Memory[6735] = 8'h01;
Memory[6734] = 8'hDE;
Memory[6733] = 8'h14;
Memory[6732] = 8'h63;
Memory[6739] = 8'h09;
Memory[6738] = 8'hC0;
Memory[6737] = 8'h00;
Memory[6736] = 8'h6F;
Memory[6743] = 8'h01;
Memory[6742] = 8'hDE;
Memory[6741] = 8'h42;
Memory[6740] = 8'h33;
Memory[6747] = 8'h01;
Memory[6746] = 8'h82;
Memory[6745] = 8'h71;
Memory[6744] = 8'hB3;
Memory[6751] = 8'h01;
Memory[6750] = 8'hD1;
Memory[6749] = 8'hF1;
Memory[6748] = 8'hB3;
Memory[6755] = 8'h00;
Memory[6754] = 8'h01;
Memory[6753] = 8'h84;
Memory[6752] = 8'h63;
Memory[6759] = 8'h0D;
Memory[6758] = 8'h00;
Memory[6757] = 8'h20;
Memory[6756] = 8'h6F;
Memory[6763] = 8'h01;
Memory[6762] = 8'h72;
Memory[6761] = 8'h71;
Memory[6760] = 8'hB3;
Memory[6767] = 8'hFF;
Memory[6766] = 8'hF0;
Memory[6765] = 8'h02;
Memory[6764] = 8'h93;
Memory[6771] = 8'h01;
Memory[6770] = 8'hD2;
Memory[6769] = 8'hC2;
Memory[6768] = 8'hB3;
Memory[6775] = 8'h00;
Memory[6774] = 8'h51;
Memory[6773] = 8'hF1;
Memory[6772] = 8'hB3;
Memory[6779] = 8'h02;
Memory[6778] = 8'h01;
Memory[6777] = 8'h94;
Memory[6776] = 8'h63;
Memory[6783] = 8'hFF;
Memory[6782] = 8'hF2;
Memory[6781] = 8'h71;
Memory[6780] = 8'h93;
Memory[6787] = 8'h01;
Memory[6786] = 8'hD1;
Memory[6785] = 8'hF1;
Memory[6784] = 8'hB3;
Memory[6791] = 8'h00;
Memory[6790] = 8'h01;
Memory[6789] = 8'h94;
Memory[6788] = 8'h63;
Memory[6795] = 8'h2C;
Memory[6794] = 8'h40;
Memory[6793] = 8'h00;
Memory[6792] = 8'h6F;
Memory[6799] = 8'h40;
Memory[6798] = 8'h01;
Memory[6797] = 8'hF2;
Memory[6796] = 8'h13;
Memory[6803] = 8'h02;
Memory[6802] = 8'h02;
Memory[6801] = 8'h10;
Memory[6800] = 8'h63;
Memory[6807] = 8'h01;
Memory[6806] = 8'h01;
Memory[6805] = 8'hF2;
Memory[6804] = 8'h13;
Memory[6811] = 8'h02;
Memory[6810] = 8'h02;
Memory[6809] = 8'h12;
Memory[6808] = 8'h63;
Memory[6815] = 8'h2C;
Memory[6814] = 8'h40;
Memory[6813] = 8'h00;
Memory[6812] = 8'h6F;
Memory[6819] = 8'h03;
Memory[6818] = 8'h20;
Memory[6817] = 8'h01;
Memory[6816] = 8'h13;
Memory[6823] = 8'h00;
Memory[6822] = 8'h0E;
Memory[6821] = 8'h8E;
Memory[6820] = 8'h13;
Memory[6827] = 8'h4A;
Memory[6826] = 8'h10;
Memory[6825] = 8'h10;
Memory[6824] = 8'h6F;
Memory[6831] = 8'h00;
Memory[6830] = 8'h0B;
Memory[6829] = 8'h2A;
Memory[6828] = 8'h23;
Memory[6835] = 8'h03;
Memory[6834] = 8'h00;
Memory[6833] = 8'h01;
Memory[6832] = 8'h13;
Memory[6839] = 8'h00;
Memory[6838] = 8'h0E;
Memory[6837] = 8'h8E;
Memory[6836] = 8'h13;
Memory[6843] = 8'h35;
Memory[6842] = 8'hD0;
Memory[6841] = 8'h10;
Memory[6840] = 8'h6F;
Memory[6847] = 8'h03;
Memory[6846] = 8'h10;
Memory[6845] = 8'h01;
Memory[6844] = 8'h13;
Memory[6851] = 8'h00;
Memory[6850] = 8'h0E;
Memory[6849] = 8'h8E;
Memory[6848] = 8'h13;
Memory[6855] = 8'h40;
Memory[6854] = 8'hD0;
Memory[6853] = 8'h10;
Memory[6852] = 8'h6F;
Memory[6859] = 8'h02;
Memory[6858] = 8'hF0;
Memory[6857] = 8'h01;
Memory[6856] = 8'h13;
Memory[6863] = 8'h20;
Memory[6862] = 8'h8B;
Memory[6861] = 8'h21;
Memory[6860] = 8'h83;
Memory[6867] = 8'h20;
Memory[6866] = 8'hCB;
Memory[6865] = 8'h22;
Memory[6864] = 8'h03;
Memory[6871] = 8'h01;
Memory[6870] = 8'hA0;
Memory[6869] = 8'h02;
Memory[6868] = 8'h93;
Memory[6875] = 8'h00;
Memory[6874] = 8'h3B;
Memory[6873] = 8'h20;
Memory[6872] = 8'h23;
Memory[6879] = 8'h00;
Memory[6878] = 8'h4B;
Memory[6877] = 8'h22;
Memory[6876] = 8'h23;
Memory[6883] = 8'h00;
Memory[6882] = 8'h5B;
Memory[6881] = 8'h24;
Memory[6880] = 8'h23;
Memory[6887] = 8'h01;
Memory[6886] = 8'hDE;
Memory[6885] = 8'h14;
Memory[6884] = 8'h63;
Memory[6891] = 8'h09;
Memory[6890] = 8'hC0;
Memory[6889] = 8'h00;
Memory[6888] = 8'h6F;
Memory[6895] = 8'h01;
Memory[6894] = 8'hDE;
Memory[6893] = 8'h42;
Memory[6892] = 8'h33;
Memory[6899] = 8'h01;
Memory[6898] = 8'h82;
Memory[6897] = 8'h71;
Memory[6896] = 8'hB3;
Memory[6903] = 8'h01;
Memory[6902] = 8'hD1;
Memory[6901] = 8'hF1;
Memory[6900] = 8'hB3;
Memory[6907] = 8'h00;
Memory[6906] = 8'h01;
Memory[6905] = 8'h84;
Memory[6904] = 8'h63;
Memory[6911] = 8'h0D;
Memory[6910] = 8'h00;
Memory[6909] = 8'h20;
Memory[6908] = 8'h6F;
Memory[6915] = 8'h01;
Memory[6914] = 8'h72;
Memory[6913] = 8'h71;
Memory[6912] = 8'hB3;
Memory[6919] = 8'hFF;
Memory[6918] = 8'hF0;
Memory[6917] = 8'h02;
Memory[6916] = 8'h93;
Memory[6923] = 8'h01;
Memory[6922] = 8'hD2;
Memory[6921] = 8'hC2;
Memory[6920] = 8'hB3;
Memory[6927] = 8'h00;
Memory[6926] = 8'h51;
Memory[6925] = 8'hF1;
Memory[6924] = 8'hB3;
Memory[6931] = 8'h02;
Memory[6930] = 8'h01;
Memory[6929] = 8'h94;
Memory[6928] = 8'h63;
Memory[6935] = 8'hFF;
Memory[6934] = 8'hF2;
Memory[6933] = 8'h71;
Memory[6932] = 8'h93;
Memory[6939] = 8'h01;
Memory[6938] = 8'hD1;
Memory[6937] = 8'hF1;
Memory[6936] = 8'hB3;
Memory[6943] = 8'h00;
Memory[6942] = 8'h01;
Memory[6941] = 8'h94;
Memory[6940] = 8'h63;
Memory[6947] = 8'h2C;
Memory[6946] = 8'h40;
Memory[6945] = 8'h00;
Memory[6944] = 8'h6F;
Memory[6951] = 8'h01;
Memory[6950] = 8'h01;
Memory[6949] = 8'hF2;
Memory[6948] = 8'h13;
Memory[6955] = 8'h00;
Memory[6954] = 8'h02;
Memory[6953] = 8'h1E;
Memory[6952] = 8'h63;
Memory[6959] = 8'h00;
Memory[6958] = 8'h41;
Memory[6957] = 8'hF2;
Memory[6956] = 8'h13;
Memory[6963] = 8'h02;
Memory[6962] = 8'h02;
Memory[6961] = 8'h10;
Memory[6960] = 8'h63;
Memory[6967] = 8'h2C;
Memory[6966] = 8'h40;
Memory[6965] = 8'h00;
Memory[6964] = 8'h6F;
Memory[6971] = 8'h03;
Memory[6970] = 8'h20;
Memory[6969] = 8'h01;
Memory[6968] = 8'h13;
Memory[6975] = 8'h00;
Memory[6974] = 8'h0E;
Memory[6973] = 8'h8E;
Memory[6972] = 8'h13;
Memory[6979] = 8'h4A;
Memory[6978] = 8'h10;
Memory[6977] = 8'h10;
Memory[6976] = 8'h6F;
Memory[6983] = 8'h03;
Memory[6982] = 8'h00;
Memory[6981] = 8'h01;
Memory[6980] = 8'h13;
Memory[6987] = 8'h00;
Memory[6986] = 8'h0E;
Memory[6985] = 8'h8E;
Memory[6984] = 8'h13;
Memory[6991] = 8'h35;
Memory[6990] = 8'hD0;
Memory[6989] = 8'h10;
Memory[6988] = 8'h6F;
Memory[6995] = 8'h03;
Memory[6994] = 8'h20;
Memory[6993] = 8'h01;
Memory[6992] = 8'h13;
Memory[6999] = 8'h00;
Memory[6998] = 8'h0E;
Memory[6997] = 8'h8E;
Memory[6996] = 8'h13;
Memory[7003] = 8'h4A;
Memory[7002] = 8'h10;
Memory[7001] = 8'h10;
Memory[7000] = 8'h6F;
Memory[7007] = 8'h03;
Memory[7006] = 8'h00;
Memory[7005] = 8'h01;
Memory[7004] = 8'h13;
Memory[7011] = 8'h20;
Memory[7010] = 8'h0B;
Memory[7009] = 8'h21;
Memory[7008] = 8'h83;
Memory[7015] = 8'h20;
Memory[7014] = 8'h4B;
Memory[7013] = 8'h22;
Memory[7012] = 8'h03;
Memory[7019] = 8'h01;
Memory[7018] = 8'hA0;
Memory[7017] = 8'h02;
Memory[7016] = 8'h93;
Memory[7023] = 8'h00;
Memory[7022] = 8'h3B;
Memory[7021] = 8'h20;
Memory[7020] = 8'h23;
Memory[7027] = 8'h00;
Memory[7026] = 8'h4B;
Memory[7025] = 8'h22;
Memory[7024] = 8'h23;
Memory[7031] = 8'h00;
Memory[7030] = 8'h5B;
Memory[7029] = 8'h24;
Memory[7028] = 8'h23;
Memory[7035] = 8'h01;
Memory[7034] = 8'hDE;
Memory[7033] = 8'h14;
Memory[7032] = 8'h63;
Memory[7039] = 8'h09;
Memory[7038] = 8'hC0;
Memory[7037] = 8'h00;
Memory[7036] = 8'h6F;
Memory[7043] = 8'h01;
Memory[7042] = 8'hDE;
Memory[7041] = 8'h42;
Memory[7040] = 8'h33;
Memory[7047] = 8'h01;
Memory[7046] = 8'h82;
Memory[7045] = 8'h71;
Memory[7044] = 8'hB3;
Memory[7051] = 8'h01;
Memory[7050] = 8'hD1;
Memory[7049] = 8'hF1;
Memory[7048] = 8'hB3;
Memory[7055] = 8'h00;
Memory[7054] = 8'h01;
Memory[7053] = 8'h84;
Memory[7052] = 8'h63;
Memory[7059] = 8'h0D;
Memory[7058] = 8'h00;
Memory[7057] = 8'h20;
Memory[7056] = 8'h6F;
Memory[7063] = 8'h01;
Memory[7062] = 8'h72;
Memory[7061] = 8'h71;
Memory[7060] = 8'hB3;
Memory[7067] = 8'hFF;
Memory[7066] = 8'hF0;
Memory[7065] = 8'h02;
Memory[7064] = 8'h93;
Memory[7071] = 8'h01;
Memory[7070] = 8'hD2;
Memory[7069] = 8'hC2;
Memory[7068] = 8'hB3;
Memory[7075] = 8'h00;
Memory[7074] = 8'h51;
Memory[7073] = 8'hF1;
Memory[7072] = 8'hB3;
Memory[7079] = 8'h02;
Memory[7078] = 8'h01;
Memory[7077] = 8'h98;
Memory[7076] = 8'h63;
Memory[7083] = 8'hFF;
Memory[7082] = 8'hF2;
Memory[7081] = 8'h71;
Memory[7080] = 8'h93;
Memory[7087] = 8'h01;
Memory[7086] = 8'hD1;
Memory[7085] = 8'hF1;
Memory[7084] = 8'hB3;
Memory[7091] = 8'h00;
Memory[7090] = 8'h01;
Memory[7089] = 8'h94;
Memory[7088] = 8'h63;
Memory[7095] = 8'h2C;
Memory[7094] = 8'h40;
Memory[7093] = 8'h00;
Memory[7092] = 8'h6F;
Memory[7099] = 8'h40;
Memory[7098] = 8'h01;
Memory[7097] = 8'hF2;
Memory[7096] = 8'h13;
Memory[7103] = 8'h02;
Memory[7102] = 8'h02;
Memory[7101] = 8'h12;
Memory[7100] = 8'h63;
Memory[7107] = 8'h01;
Memory[7106] = 8'h01;
Memory[7105] = 8'hF2;
Memory[7104] = 8'h13;
Memory[7111] = 8'h02;
Memory[7110] = 8'h02;
Memory[7109] = 8'h14;
Memory[7108] = 8'h63;
Memory[7115] = 8'h00;
Memory[7114] = 8'h41;
Memory[7113] = 8'hF2;
Memory[7112] = 8'h13;
Memory[7119] = 8'h02;
Memory[7118] = 8'h02;
Memory[7117] = 8'h16;
Memory[7116] = 8'h63;
Memory[7123] = 8'h2C;
Memory[7122] = 8'h40;
Memory[7121] = 8'h00;
Memory[7120] = 8'h6F;
Memory[7127] = 8'h03;
Memory[7126] = 8'h20;
Memory[7125] = 8'h01;
Memory[7124] = 8'h13;
Memory[7131] = 8'h00;
Memory[7130] = 8'h0E;
Memory[7129] = 8'h8E;
Memory[7128] = 8'h13;
Memory[7135] = 8'h4A;
Memory[7134] = 8'h10;
Memory[7133] = 8'h10;
Memory[7132] = 8'h6F;
Memory[7139] = 8'h02;
Memory[7138] = 8'hF0;
Memory[7137] = 8'h01;
Memory[7136] = 8'h13;
Memory[7143] = 8'h00;
Memory[7142] = 8'h0E;
Memory[7141] = 8'h8E;
Memory[7140] = 8'h13;
Memory[7147] = 8'h2C;
Memory[7146] = 8'h90;
Memory[7145] = 8'h10;
Memory[7144] = 8'h6F;
Memory[7151] = 8'h02;
Memory[7150] = 8'hE0;
Memory[7149] = 8'h01;
Memory[7148] = 8'h13;
Memory[7155] = 8'h00;
Memory[7154] = 8'h0E;
Memory[7153] = 8'h8E;
Memory[7152] = 8'h13;
Memory[7159] = 8'h23;
Memory[7158] = 8'h10;
Memory[7157] = 8'h10;
Memory[7156] = 8'h6F;
Memory[7163] = 8'h02;
Memory[7162] = 8'hB0;
Memory[7161] = 8'h01;
Memory[7160] = 8'h13;
Memory[7167] = 8'h00;
Memory[7166] = 8'h0E;
Memory[7165] = 8'h8E;
Memory[7164] = 8'h13;
Memory[7171] = 8'h08;
Memory[7170] = 8'h0B;
Memory[7169] = 8'h2E;
Memory[7168] = 8'h23;
Memory[7175] = 8'h05;
Memory[7174] = 8'hFB;
Memory[7173] = 8'h28;
Memory[7172] = 8'h23;
Memory[7179] = 8'h1E;
Memory[7178] = 8'h50;
Memory[7177] = 8'h10;
Memory[7176] = 8'h6F;
Memory[7183] = 8'h03;
Memory[7182] = 8'h10;
Memory[7181] = 8'h01;
Memory[7180] = 8'h13;
Memory[7187] = 8'h21;
Memory[7186] = 8'h0B;
Memory[7185] = 8'h21;
Memory[7184] = 8'h83;
Memory[7191] = 8'h21;
Memory[7190] = 8'h4B;
Memory[7189] = 8'h22;
Memory[7188] = 8'h03;
Memory[7195] = 8'h01;
Memory[7194] = 8'h90;
Memory[7193] = 8'h02;
Memory[7192] = 8'h93;
Memory[7199] = 8'h00;
Memory[7198] = 8'h3B;
Memory[7197] = 8'h20;
Memory[7196] = 8'h23;
Memory[7203] = 8'h00;
Memory[7202] = 8'h4B;
Memory[7201] = 8'h22;
Memory[7200] = 8'h23;
Memory[7207] = 8'h00;
Memory[7206] = 8'h5B;
Memory[7205] = 8'h24;
Memory[7204] = 8'h23;
Memory[7211] = 8'h01;
Memory[7210] = 8'hDE;
Memory[7209] = 8'h14;
Memory[7208] = 8'h63;
Memory[7215] = 8'h09;
Memory[7214] = 8'hC0;
Memory[7213] = 8'h00;
Memory[7212] = 8'h6F;
Memory[7219] = 8'h01;
Memory[7218] = 8'hDE;
Memory[7217] = 8'h42;
Memory[7216] = 8'h33;
Memory[7223] = 8'h01;
Memory[7222] = 8'h82;
Memory[7221] = 8'h71;
Memory[7220] = 8'hB3;
Memory[7227] = 8'h01;
Memory[7226] = 8'hD1;
Memory[7225] = 8'hF1;
Memory[7224] = 8'hB3;
Memory[7231] = 8'h00;
Memory[7230] = 8'h01;
Memory[7229] = 8'h84;
Memory[7228] = 8'h63;
Memory[7235] = 8'h0D;
Memory[7234] = 8'h00;
Memory[7233] = 8'h20;
Memory[7232] = 8'h6F;
Memory[7239] = 8'h01;
Memory[7238] = 8'h72;
Memory[7237] = 8'h71;
Memory[7236] = 8'hB3;
Memory[7243] = 8'hFF;
Memory[7242] = 8'hF0;
Memory[7241] = 8'h02;
Memory[7240] = 8'h93;
Memory[7247] = 8'h01;
Memory[7246] = 8'hD2;
Memory[7245] = 8'hC2;
Memory[7244] = 8'hB3;
Memory[7251] = 8'h00;
Memory[7250] = 8'h51;
Memory[7249] = 8'hF1;
Memory[7248] = 8'hB3;
Memory[7255] = 8'h02;
Memory[7254] = 8'h01;
Memory[7253] = 8'h94;
Memory[7252] = 8'h63;
Memory[7259] = 8'hFF;
Memory[7258] = 8'hF2;
Memory[7257] = 8'h71;
Memory[7256] = 8'h93;
Memory[7263] = 8'h01;
Memory[7262] = 8'hD1;
Memory[7261] = 8'hF1;
Memory[7260] = 8'hB3;
Memory[7267] = 8'h00;
Memory[7266] = 8'h01;
Memory[7265] = 8'h94;
Memory[7264] = 8'h63;
Memory[7271] = 8'h2C;
Memory[7270] = 8'h40;
Memory[7269] = 8'h00;
Memory[7268] = 8'h6F;
Memory[7275] = 8'h40;
Memory[7274] = 8'h01;
Memory[7273] = 8'hF2;
Memory[7272] = 8'h13;
Memory[7279] = 8'h00;
Memory[7278] = 8'h02;
Memory[7277] = 8'h1E;
Memory[7276] = 8'h63;
Memory[7283] = 8'h00;
Memory[7282] = 8'h41;
Memory[7281] = 8'hF2;
Memory[7280] = 8'h13;
Memory[7287] = 8'h02;
Memory[7286] = 8'h02;
Memory[7285] = 8'h10;
Memory[7284] = 8'h63;
Memory[7291] = 8'h2C;
Memory[7290] = 8'h40;
Memory[7289] = 8'h00;
Memory[7288] = 8'h6F;
Memory[7295] = 8'h03;
Memory[7294] = 8'h20;
Memory[7293] = 8'h01;
Memory[7292] = 8'h13;
Memory[7299] = 8'h00;
Memory[7298] = 8'h0E;
Memory[7297] = 8'h8E;
Memory[7296] = 8'h13;
Memory[7303] = 8'h4A;
Memory[7302] = 8'h10;
Memory[7301] = 8'h10;
Memory[7300] = 8'h6F;
Memory[7307] = 8'h02;
Memory[7306] = 8'hE0;
Memory[7305] = 8'h01;
Memory[7304] = 8'h13;
Memory[7311] = 8'h00;
Memory[7310] = 8'h0E;
Memory[7309] = 8'h8E;
Memory[7308] = 8'h13;
Memory[7315] = 8'h23;
Memory[7314] = 8'h10;
Memory[7313] = 8'h10;
Memory[7312] = 8'h6F;
Memory[7319] = 8'h00;
Memory[7318] = 8'h80;
Memory[7317] = 8'h01;
Memory[7316] = 8'h13;
Memory[7323] = 8'h00;
Memory[7322] = 8'h0E;
Memory[7321] = 8'h8E;
Memory[7320] = 8'h13;
Memory[7327] = 8'h6A;
Memory[7326] = 8'h80;
Memory[7325] = 8'h00;
Memory[7324] = 8'h6F;
Memory[7331] = 8'h03;
Memory[7330] = 8'h20;
Memory[7329] = 8'h01;
Memory[7328] = 8'h13;
Memory[7335] = 8'h23;
Memory[7334] = 8'h0B;
Memory[7333] = 8'h21;
Memory[7332] = 8'h83;
Memory[7339] = 8'h23;
Memory[7338] = 8'h4B;
Memory[7337] = 8'h22;
Memory[7336] = 8'h03;
Memory[7343] = 8'h01;
Memory[7342] = 8'h80;
Memory[7341] = 8'h02;
Memory[7340] = 8'h93;
Memory[7347] = 8'h00;
Memory[7346] = 8'h3B;
Memory[7345] = 8'h20;
Memory[7344] = 8'h23;
Memory[7351] = 8'h00;
Memory[7350] = 8'h4B;
Memory[7349] = 8'h22;
Memory[7348] = 8'h23;
Memory[7355] = 8'h00;
Memory[7354] = 8'h5B;
Memory[7353] = 8'h24;
Memory[7352] = 8'h23;
Memory[7359] = 8'h01;
Memory[7358] = 8'hDE;
Memory[7357] = 8'h14;
Memory[7356] = 8'h63;
Memory[7363] = 8'h09;
Memory[7362] = 8'hC0;
Memory[7361] = 8'h00;
Memory[7360] = 8'h6F;
Memory[7367] = 8'h01;
Memory[7366] = 8'hDE;
Memory[7365] = 8'h42;
Memory[7364] = 8'h33;
Memory[7371] = 8'h01;
Memory[7370] = 8'h82;
Memory[7369] = 8'h71;
Memory[7368] = 8'hB3;
Memory[7375] = 8'h01;
Memory[7374] = 8'hD1;
Memory[7373] = 8'hF1;
Memory[7372] = 8'hB3;
Memory[7379] = 8'h00;
Memory[7378] = 8'h01;
Memory[7377] = 8'h84;
Memory[7376] = 8'h63;
Memory[7383] = 8'h0D;
Memory[7382] = 8'h00;
Memory[7381] = 8'h20;
Memory[7380] = 8'h6F;
Memory[7387] = 8'hFF;
Memory[7386] = 8'hF2;
Memory[7385] = 8'h71;
Memory[7384] = 8'h93;
Memory[7391] = 8'h01;
Memory[7390] = 8'hD1;
Memory[7389] = 8'hF1;
Memory[7388] = 8'hB3;
Memory[7395] = 8'h00;
Memory[7394] = 8'h01;
Memory[7393] = 8'h94;
Memory[7392] = 8'h63;
Memory[7399] = 8'h2C;
Memory[7398] = 8'h40;
Memory[7397] = 8'h00;
Memory[7396] = 8'h6F;
Memory[7403] = 8'h02;
Memory[7402] = 8'hB0;
Memory[7401] = 8'h01;
Memory[7400] = 8'h13;
Memory[7407] = 8'h00;
Memory[7406] = 8'h0E;
Memory[7405] = 8'h8E;
Memory[7404] = 8'h13;
Memory[7411] = 8'h05;
Memory[7410] = 8'h0B;
Memory[7409] = 8'h21;
Memory[7408] = 8'h83;
Memory[7415] = 8'h09;
Memory[7414] = 8'hCB;
Memory[7413] = 8'h22;
Memory[7412] = 8'h03;
Memory[7419] = 8'h40;
Memory[7418] = 8'h32;
Memory[7417] = 8'h01;
Memory[7416] = 8'hB3;
Memory[7423] = 8'h40;
Memory[7422] = 8'h3F;
Memory[7421] = 8'h81;
Memory[7420] = 8'hB3;
Memory[7427] = 8'h04;
Memory[7426] = 8'h3B;
Memory[7425] = 8'h28;
Memory[7424] = 8'h23;
Memory[7431] = 8'h1E;
Memory[7430] = 8'h50;
Memory[7429] = 8'h10;
Memory[7428] = 8'h6F;
Memory[7435] = 8'h03;
Memory[7434] = 8'h40;
Memory[7433] = 8'h01;
Memory[7432] = 8'h13;
Memory[7439] = 8'h22;
Memory[7438] = 8'h8B;
Memory[7437] = 8'h21;
Memory[7436] = 8'h83;
Memory[7443] = 8'h22;
Memory[7442] = 8'hCB;
Memory[7441] = 8'h22;
Memory[7440] = 8'h03;
Memory[7447] = 8'h00;
Memory[7446] = 8'hC0;
Memory[7445] = 8'h02;
Memory[7444] = 8'h93;
Memory[7451] = 8'h00;
Memory[7450] = 8'h3B;
Memory[7449] = 8'h20;
Memory[7448] = 8'h23;
Memory[7455] = 8'h00;
Memory[7454] = 8'h4B;
Memory[7453] = 8'h22;
Memory[7452] = 8'h23;
Memory[7459] = 8'h00;
Memory[7458] = 8'h5B;
Memory[7457] = 8'h24;
Memory[7456] = 8'h23;
Memory[7463] = 8'h01;
Memory[7462] = 8'hDE;
Memory[7461] = 8'h14;
Memory[7460] = 8'h63;
Memory[7467] = 8'h09;
Memory[7466] = 8'hC0;
Memory[7465] = 8'h00;
Memory[7464] = 8'h6F;
Memory[7471] = 8'h01;
Memory[7470] = 8'hDE;
Memory[7469] = 8'h42;
Memory[7468] = 8'h33;
Memory[7475] = 8'h01;
Memory[7474] = 8'h82;
Memory[7473] = 8'h71;
Memory[7472] = 8'hB3;
Memory[7479] = 8'h01;
Memory[7478] = 8'hD1;
Memory[7477] = 8'hF1;
Memory[7476] = 8'hB3;
Memory[7483] = 8'h00;
Memory[7482] = 8'h01;
Memory[7481] = 8'h84;
Memory[7480] = 8'h63;
Memory[7487] = 8'h0D;
Memory[7486] = 8'h00;
Memory[7485] = 8'h20;
Memory[7484] = 8'h6F;
Memory[7491] = 8'hFF;
Memory[7490] = 8'hF2;
Memory[7489] = 8'h71;
Memory[7488] = 8'h93;
Memory[7495] = 8'h01;
Memory[7494] = 8'hD1;
Memory[7493] = 8'hF1;
Memory[7492] = 8'hB3;
Memory[7499] = 8'h00;
Memory[7498] = 8'h01;
Memory[7497] = 8'h94;
Memory[7496] = 8'h63;
Memory[7503] = 8'h2C;
Memory[7502] = 8'h40;
Memory[7501] = 8'h00;
Memory[7500] = 8'h6F;
Memory[7507] = 8'h03;
Memory[7506] = 8'h60;
Memory[7505] = 8'h01;
Memory[7504] = 8'h13;
Memory[7511] = 8'h00;
Memory[7510] = 8'h0E;
Memory[7509] = 8'h8E;
Memory[7508] = 8'h13;
Memory[7515] = 8'h55;
Memory[7514] = 8'hD0;
Memory[7513] = 8'h10;
Memory[7512] = 8'h6F;
Memory[7519] = 8'h03;
Memory[7518] = 8'h60;
Memory[7517] = 8'h01;
Memory[7516] = 8'h13;
Memory[7523] = 8'h21;
Memory[7522] = 8'h8B;
Memory[7521] = 8'h21;
Memory[7520] = 8'h83;
Memory[7527] = 8'h21;
Memory[7526] = 8'hCB;
Memory[7525] = 8'h22;
Memory[7524] = 8'h03;
Memory[7531] = 8'h01;
Memory[7530] = 8'hB0;
Memory[7529] = 8'h02;
Memory[7528] = 8'h93;
Memory[7535] = 8'h00;
Memory[7534] = 8'h3B;
Memory[7533] = 8'h20;
Memory[7532] = 8'h23;
Memory[7539] = 8'h00;
Memory[7538] = 8'h4B;
Memory[7537] = 8'h22;
Memory[7536] = 8'h23;
Memory[7543] = 8'h00;
Memory[7542] = 8'h5B;
Memory[7541] = 8'h24;
Memory[7540] = 8'h23;
Memory[7547] = 8'h01;
Memory[7546] = 8'hDE;
Memory[7545] = 8'h14;
Memory[7544] = 8'h63;
Memory[7551] = 8'h09;
Memory[7550] = 8'hC0;
Memory[7549] = 8'h00;
Memory[7548] = 8'h6F;
Memory[7555] = 8'h01;
Memory[7554] = 8'hDE;
Memory[7553] = 8'h42;
Memory[7552] = 8'h33;
Memory[7559] = 8'h01;
Memory[7558] = 8'h82;
Memory[7557] = 8'h71;
Memory[7556] = 8'hB3;
Memory[7563] = 8'h01;
Memory[7562] = 8'hD1;
Memory[7561] = 8'hF1;
Memory[7560] = 8'hB3;
Memory[7567] = 8'h00;
Memory[7566] = 8'h01;
Memory[7565] = 8'h84;
Memory[7564] = 8'h63;
Memory[7571] = 8'h0D;
Memory[7570] = 8'h00;
Memory[7569] = 8'h20;
Memory[7568] = 8'h6F;
Memory[7575] = 8'hFF;
Memory[7574] = 8'hF2;
Memory[7573] = 8'h71;
Memory[7572] = 8'h93;
Memory[7579] = 8'h01;
Memory[7578] = 8'hD1;
Memory[7577] = 8'hF1;
Memory[7576] = 8'hB3;
Memory[7583] = 8'h00;
Memory[7582] = 8'h01;
Memory[7581] = 8'h94;
Memory[7580] = 8'h63;
Memory[7587] = 8'h2C;
Memory[7586] = 8'h40;
Memory[7585] = 8'h00;
Memory[7584] = 8'h6F;
Memory[7591] = 8'h03;
Memory[7590] = 8'h70;
Memory[7589] = 8'h01;
Memory[7588] = 8'h13;
Memory[7595] = 8'h00;
Memory[7594] = 8'h0E;
Memory[7593] = 8'h8E;
Memory[7592] = 8'h13;
Memory[7599] = 8'h5B;
Memory[7598] = 8'h10;
Memory[7597] = 8'h10;
Memory[7596] = 8'h6F;
Memory[7603] = 8'h03;
Memory[7602] = 8'h70;
Memory[7601] = 8'h01;
Memory[7600] = 8'h13;
Memory[7607] = 8'h24;
Memory[7606] = 8'h0B;
Memory[7605] = 8'h21;
Memory[7604] = 8'h83;
Memory[7611] = 8'h07;
Memory[7610] = 8'h4B;
Memory[7609] = 8'h23;
Memory[7608] = 8'h83;
Memory[7615] = 8'h06;
Memory[7614] = 8'h40;
Memory[7613] = 8'h02;
Memory[7612] = 8'h93;
Memory[7619] = 8'h03;
Memory[7618] = 8'hB2;
Memory[7617] = 8'h82;
Memory[7616] = 8'hB3;
Memory[7623] = 8'h02;
Memory[7622] = 8'h53;
Memory[7621] = 8'hC2;
Memory[7620] = 8'h33;
Memory[7627] = 8'h00;
Memory[7626] = 8'hA0;
Memory[7625] = 8'h02;
Memory[7624] = 8'h93;
Memory[7631] = 8'h02;
Memory[7630] = 8'h52;
Memory[7629] = 8'h62;
Memory[7628] = 8'h33;
Memory[7635] = 8'h00;
Memory[7634] = 8'h82;
Memory[7633] = 8'h12;
Memory[7632] = 8'h13;
Memory[7639] = 8'h03;
Memory[7638] = 8'hB2;
Memory[7637] = 8'h82;
Memory[7636] = 8'hB3;
Memory[7643] = 8'h02;
Memory[7642] = 8'h53;
Memory[7641] = 8'hC3;
Memory[7640] = 8'h33;
Memory[7647] = 8'h00;
Memory[7646] = 8'hA0;
Memory[7645] = 8'h02;
Memory[7644] = 8'h93;
Memory[7651] = 8'h02;
Memory[7650] = 8'h53;
Memory[7649] = 8'h63;
Memory[7648] = 8'h33;
Memory[7655] = 8'h00;
Memory[7654] = 8'h62;
Memory[7653] = 8'h02;
Memory[7652] = 8'h33;
Memory[7659] = 8'h00;
Memory[7658] = 8'h41;
Memory[7657] = 8'h81;
Memory[7656] = 8'hB3;
Memory[7663] = 8'h00;
Memory[7662] = 8'h3B;
Memory[7661] = 8'h20;
Memory[7660] = 8'h23;
Memory[7667] = 8'h24;
Memory[7666] = 8'h4B;
Memory[7665] = 8'h21;
Memory[7664] = 8'h83;
Memory[7671] = 8'h03;
Memory[7670] = 8'hB3;
Memory[7669] = 8'hC2;
Memory[7668] = 8'h33;
Memory[7675] = 8'h02;
Memory[7674] = 8'h52;
Memory[7673] = 8'h62;
Memory[7672] = 8'h33;
Memory[7679] = 8'h00;
Memory[7678] = 8'h82;
Memory[7677] = 8'h12;
Memory[7676] = 8'h13;
Memory[7683] = 8'h06;
Memory[7682] = 8'h40;
Memory[7681] = 8'h02;
Memory[7680] = 8'h93;
Memory[7687] = 8'h02;
Memory[7686] = 8'h53;
Memory[7685] = 8'hC3;
Memory[7684] = 8'h33;
Memory[7691] = 8'h00;
Memory[7690] = 8'hA0;
Memory[7689] = 8'h02;
Memory[7688] = 8'h93;
Memory[7695] = 8'h02;
Memory[7694] = 8'h53;
Memory[7693] = 8'h63;
Memory[7692] = 8'h33;
Memory[7699] = 8'h00;
Memory[7698] = 8'h62;
Memory[7697] = 8'h02;
Memory[7696] = 8'h33;
Memory[7703] = 8'h00;
Memory[7702] = 8'h82;
Memory[7701] = 8'h12;
Memory[7700] = 8'h13;
Memory[7707] = 8'h02;
Memory[7706] = 8'h53;
Memory[7705] = 8'hC3;
Memory[7704] = 8'h33;
Memory[7711] = 8'h02;
Memory[7710] = 8'h53;
Memory[7709] = 8'h63;
Memory[7708] = 8'h33;
Memory[7715] = 8'h00;
Memory[7714] = 8'h62;
Memory[7713] = 8'h02;
Memory[7712] = 8'h33;
Memory[7719] = 8'h00;
Memory[7718] = 8'h82;
Memory[7717] = 8'h12;
Memory[7716] = 8'h13;
Memory[7723] = 8'h02;
Memory[7722] = 8'h53;
Memory[7721] = 8'hE3;
Memory[7720] = 8'h33;
Memory[7727] = 8'h00;
Memory[7726] = 8'h62;
Memory[7725] = 8'h02;
Memory[7724] = 8'h33;
Memory[7731] = 8'h00;
Memory[7730] = 8'h4B;
Memory[7729] = 8'h22;
Memory[7728] = 8'h23;
Memory[7735] = 8'h01;
Memory[7734] = 8'hDE;
Memory[7733] = 8'h14;
Memory[7732] = 8'h63;
Memory[7739] = 8'h09;
Memory[7738] = 8'hC0;
Memory[7737] = 8'h00;
Memory[7736] = 8'h6F;
Memory[7743] = 8'h01;
Memory[7742] = 8'hDE;
Memory[7741] = 8'h42;
Memory[7740] = 8'h33;
Memory[7747] = 8'h01;
Memory[7746] = 8'h82;
Memory[7745] = 8'h71;
Memory[7744] = 8'hB3;
Memory[7751] = 8'h01;
Memory[7750] = 8'hD1;
Memory[7749] = 8'hF1;
Memory[7748] = 8'hB3;
Memory[7755] = 8'h00;
Memory[7754] = 8'h01;
Memory[7753] = 8'h84;
Memory[7752] = 8'h63;
Memory[7759] = 8'h0D;
Memory[7758] = 8'h00;
Memory[7757] = 8'h20;
Memory[7756] = 8'h6F;
Memory[7763] = 8'hFF;
Memory[7762] = 8'hF2;
Memory[7761] = 8'h71;
Memory[7760] = 8'h93;
Memory[7767] = 8'h01;
Memory[7766] = 8'hD1;
Memory[7765] = 8'hF1;
Memory[7764] = 8'hB3;
Memory[7771] = 8'h00;
Memory[7770] = 8'h01;
Memory[7769] = 8'h94;
Memory[7768] = 8'h63;
Memory[7775] = 8'h2C;
Memory[7774] = 8'h40;
Memory[7773] = 8'h00;
Memory[7772] = 8'h6F;
Memory[7779] = 8'h00;
Memory[7778] = 8'h90;
Memory[7777] = 8'h01;
Memory[7776] = 8'h13;
Memory[7783] = 8'h00;
Memory[7782] = 8'h0E;
Memory[7781] = 8'h8E;
Memory[7780] = 8'h13;
Memory[7787] = 8'h71;
Memory[7786] = 8'h80;
Memory[7785] = 8'h00;
Memory[7784] = 8'h6F;
Memory[7791] = 8'hFF;
Memory[7790] = 8'hFF;
Memory[7789] = 8'hFF;
Memory[7788] = 8'hFF;
Memory[7795] = 8'hFF;
Memory[7794] = 8'hFF;
Memory[7793] = 8'hFF;
Memory[7792] = 8'hFF;
Memory[7799] = 8'h00;
Memory[7798] = 8'h00;
Memory[7797] = 8'h00;
Memory[7796] = 8'hFF;
Memory[7803] = 8'h00;
Memory[7802] = 8'h00;
Memory[7801] = 8'h80;
Memory[7800] = 8'h80;
Memory[7807] = 8'h00;
Memory[7806] = 8'h00;
Memory[7805] = 8'h00;
Memory[7804] = 8'hAA;
Memory[7811] = 8'h00;
Memory[7810] = 8'h00;
Memory[7809] = 8'h00;
Memory[7808] = 8'h00;
Memory[7815] = 8'h00;
Memory[7814] = 8'h00;
Memory[7813] = 8'h00;
Memory[7812] = 8'h7F;
Memory[7819] = 8'h00;
Memory[7818] = 8'h00;
Memory[7817] = 8'h00;
Memory[7816] = 8'h01;
Memory[7823] = 8'h00;
Memory[7822] = 8'h00;
Memory[7821] = 8'h00;
Memory[7820] = 8'h0A;
Memory[7827] = 8'h00;
Memory[7826] = 8'h00;
Memory[7825] = 8'h00;
Memory[7824] = 8'h64;
Memory[7831] = 8'h00;
Memory[7830] = 8'h00;
Memory[7829] = 8'h03;
Memory[7828] = 8'hE8;
Memory[7835] = 8'h00;
Memory[7834] = 8'h00;
Memory[7833] = 8'h27;
Memory[7832] = 8'h10;
Memory[7839] = 8'h00;
Memory[7838] = 8'h01;
Memory[7837] = 8'h86;
Memory[7836] = 8'hA0;
Memory[7843] = 8'h00;
Memory[7842] = 8'h0F;
Memory[7841] = 8'h42;
Memory[7840] = 8'h40;
Memory[7847] = 8'h00;
Memory[7846] = 8'h4C;
Memory[7845] = 8'h4B;
Memory[7844] = 8'h40;
Memory[7851] = 8'h00;
Memory[7850] = 8'h98;
Memory[7849] = 8'h96;
Memory[7848] = 8'h80;
Memory[7855] = 8'h02;
Memory[7854] = 8'hFA;
Memory[7853] = 8'hF0;
Memory[7852] = 8'h80;
Memory[7859] = 8'h05;
Memory[7858] = 8'hF5;
Memory[7857] = 8'hE1;
Memory[7856] = 8'h00;
Memory[7863] = 8'h1D;
Memory[7862] = 8'hCD;
Memory[7861] = 8'h65;
Memory[7860] = 8'h00;
Memory[7867] = 8'h3B;
Memory[7866] = 8'h9A;
Memory[7865] = 8'hCA;
Memory[7864] = 8'h00;
Memory[7871] = 8'h00;
Memory[7870] = 8'h00;
Memory[7869] = 8'h00;
Memory[7868] = 8'h00;
Memory[7875] = 8'h00;
Memory[7874] = 8'h02;
Memory[7873] = 8'h5D;
Memory[7872] = 8'h78;
Memory[7879] = 8'h00;
Memory[7878] = 8'h00;
Memory[7877] = 8'h00;
Memory[7876] = 8'h00;
Memory[7883] = 8'h00;
Memory[7882] = 8'h00;
Memory[7881] = 8'h00;
Memory[7880] = 8'h00;
Memory[7887] = 8'h00;
Memory[7886] = 8'h00;
Memory[7885] = 8'h00;
Memory[7884] = 8'h00;
Memory[7891] = 8'h00;
Memory[7890] = 8'h00;
Memory[7889] = 8'h00;
Memory[7888] = 8'h00;
Memory[7895] = 8'h00;
Memory[7894] = 8'h00;
Memory[7893] = 8'h00;
Memory[7892] = 8'h00;
Memory[7899] = 8'h00;
Memory[7898] = 8'h00;
Memory[7897] = 8'h00;
Memory[7896] = 8'h00;
Memory[7903] = 8'h00;
Memory[7902] = 8'h00;
Memory[7901] = 8'h00;
Memory[7900] = 8'h00;
Memory[7907] = 8'h00;
Memory[7906] = 8'h00;
Memory[7905] = 8'h00;
Memory[7904] = 8'h00;
Memory[7911] = 8'h00;
Memory[7910] = 8'h00;
Memory[7909] = 8'h00;
Memory[7908] = 8'h00;
Memory[7915] = 8'h00;
Memory[7914] = 8'h00;
Memory[7913] = 8'h00;
Memory[7912] = 8'h00;
Memory[7919] = 8'h00;
Memory[7918] = 8'h00;
Memory[7917] = 8'h00;
Memory[7916] = 8'h00;
Memory[7923] = 8'h00;
Memory[7922] = 8'h00;
Memory[7921] = 8'h00;
Memory[7920] = 8'h00;
Memory[7927] = 8'h00;
Memory[7926] = 8'h00;
Memory[7925] = 8'h00;
Memory[7924] = 8'h00;
Memory[7931] = 8'h00;
Memory[7930] = 8'h00;
Memory[7929] = 8'h00;
Memory[7928] = 8'h00;
Memory[7935] = 8'h00;
Memory[7934] = 8'h00;
Memory[7933] = 8'h00;
Memory[7932] = 8'h00;
Memory[7939] = 8'h00;
Memory[7938] = 8'h00;
Memory[7937] = 8'h00;
Memory[7936] = 8'h00;
Memory[7943] = 8'h05;
Memory[7942] = 8'hF5;
Memory[7941] = 8'hE1;
Memory[7940] = 8'h00;
Memory[7947] = 8'h00;
Memory[7946] = 8'h00;
Memory[7945] = 8'h00;
Memory[7944] = 8'h00;
Memory[7951] = 8'h24;
Memory[7950] = 8'h24;
Memory[7949] = 8'h24;
Memory[7948] = 8'h11;
Memory[7955] = 8'h0E;
Memory[7954] = 8'h15;
Memory[7953] = 8'h15;
Memory[7952] = 8'h17;
Memory[7959] = 8'h0F;
Memory[7958] = 8'h1A;
Memory[7957] = 8'h0E;
Memory[7956] = 8'h19;
Memory[7963] = 8'h1D;
Memory[7962] = 8'h16;
Memory[7961] = 8'h0C;
Memory[7960] = 8'h1F;
Memory[7967] = 8'h24;
Memory[7966] = 8'h24;
Memory[7965] = 8'h24;
Memory[7964] = 8'h01;
Memory[7971] = 8'h16;
Memory[7970] = 8'h16;
Memory[7969] = 8'h11;
Memory[7968] = 8'h20;
Memory[7975] = 8'h24;
Memory[7974] = 8'h24;
Memory[7973] = 8'h01;
Memory[7972] = 8'h00;
Memory[7979] = 8'h16;
Memory[7978] = 8'h16;
Memory[7977] = 8'h11;
Memory[7976] = 8'h20;
Memory[7983] = 8'h24;
Memory[7982] = 8'h24;
Memory[7981] = 8'h05;
Memory[7980] = 8'h00;
Memory[7987] = 8'h16;
Memory[7986] = 8'h16;
Memory[7985] = 8'h11;
Memory[7984] = 8'h20;
Memory[7991] = 8'h24;
Memory[7990] = 8'h01;
Memory[7989] = 8'h00;
Memory[7988] = 8'h00;
Memory[7995] = 8'h16;
Memory[7994] = 8'h16;
Memory[7993] = 8'h11;
Memory[7992] = 8'h20;
Memory[7999] = 8'h24;
Memory[7998] = 8'h05;
Memory[7997] = 8'h00;
Memory[7996] = 8'h00;
Memory[8003] = 8'h16;
Memory[8002] = 8'h16;
Memory[8001] = 8'h11;
Memory[8000] = 8'h20;
Memory[8007] = 8'h24;
Memory[8006] = 8'h24;
Memory[8005] = 8'h24;
Memory[8004] = 8'h01;
Memory[8011] = 8'h22;
Memory[8010] = 8'h10;
Memory[8009] = 8'h11;
Memory[8008] = 8'h20;
Memory[8015] = 8'h24;
Memory[8014] = 8'h24;
Memory[8013] = 8'h24;
Memory[8012] = 8'h1B;
Memory[8019] = 8'h1C;
Memory[8018] = 8'h0A;
Memory[8017] = 8'h1A;
Memory[8016] = 8'h1C;
Memory[8023] = 8'h24;
Memory[8022] = 8'h24;
Memory[8021] = 8'h24;
Memory[8020] = 8'h1B;
Memory[8027] = 8'h0C;
Memory[8026] = 8'h17;
Memory[8025] = 8'h1A;
Memory[8024] = 8'h0E;
Memory[8031] = 8'h01;
Memory[8030] = 8'h24;
Memory[8029] = 8'h00;
Memory[8028] = 8'h00;
Memory[8035] = 8'h00;
Memory[8034] = 8'h00;
Memory[8033] = 8'h00;
Memory[8032] = 8'h00;
Memory[8039] = 8'h02;
Memory[8038] = 8'h24;
Memory[8037] = 8'h00;
Memory[8036] = 8'h00;
Memory[8043] = 8'h00;
Memory[8042] = 8'h00;
Memory[8041] = 8'h00;
Memory[8040] = 8'h00;
Memory[8047] = 8'h03;
Memory[8046] = 8'h24;
Memory[8045] = 8'h00;
Memory[8044] = 8'h00;
Memory[8051] = 8'h00;
Memory[8050] = 8'h00;
Memory[8049] = 8'h00;
Memory[8048] = 8'h00;
Memory[8055] = 8'h04;
Memory[8054] = 8'h24;
Memory[8053] = 8'h00;
Memory[8052] = 8'h00;
Memory[8059] = 8'h00;
Memory[8058] = 8'h00;
Memory[8057] = 8'h00;
Memory[8056] = 8'h00;
Memory[8063] = 8'h05;
Memory[8062] = 8'h24;
Memory[8061] = 8'h00;
Memory[8060] = 8'h00;
Memory[8067] = 8'h00;
Memory[8066] = 8'h00;
Memory[8065] = 8'h00;
Memory[8064] = 8'h00;
Memory[8071] = 8'h06;
Memory[8070] = 8'h24;
Memory[8069] = 8'h00;
Memory[8068] = 8'h00;
Memory[8075] = 8'h00;
Memory[8074] = 8'h00;
Memory[8073] = 8'h00;
Memory[8072] = 8'h00;
Memory[8079] = 8'h07;
Memory[8078] = 8'h24;
Memory[8077] = 8'h00;
Memory[8076] = 8'h00;
Memory[8083] = 8'h00;
Memory[8082] = 8'h00;
Memory[8081] = 8'h00;
Memory[8080] = 8'h00;
Memory[8087] = 8'h08;
Memory[8086] = 8'h24;
Memory[8085] = 8'h00;
Memory[8084] = 8'h00;
Memory[8091] = 8'h00;
Memory[8090] = 8'h00;
Memory[8089] = 8'h00;
Memory[8088] = 8'h00;
Memory[8095] = 8'h09;
Memory[8094] = 8'h24;
Memory[8093] = 8'h00;
Memory[8092] = 8'h00;
Memory[8099] = 8'h00;
Memory[8098] = 8'h00;
Memory[8097] = 8'h00;
Memory[8096] = 8'h00;
Memory[8103] = 8'h24;
Memory[8102] = 8'h24;
Memory[8101] = 8'h24;
Memory[8100] = 8'h24;
Memory[8107] = 8'h12;
Memory[8106] = 8'h16;
Memory[8105] = 8'h0F;
Memory[8104] = 8'h17;
Memory[8111] = 8'h24;
Memory[8110] = 8'h1A;
Memory[8109] = 8'h11;
Memory[8108] = 8'h1F;
Memory[8115] = 8'h1C;
Memory[8114] = 8'h11;
Memory[8113] = 8'h16;
Memory[8112] = 8'h16;
Memory[8119] = 8'h24;
Memory[8118] = 8'h24;
Memory[8117] = 8'h10;
Memory[8116] = 8'h0A;
Memory[8123] = 8'h16;
Memory[8122] = 8'h16;
Memory[8121] = 8'h0E;
Memory[8120] = 8'h24;
Memory[8127] = 8'h0D;
Memory[8126] = 8'h0E;
Memory[8125] = 8'h1E;
Memory[8124] = 8'h15;
Memory[8131] = 8'h17;
Memory[8130] = 8'h18;
Memory[8129] = 8'h0E;
Memory[8128] = 8'h0D;
Memory[8135] = 8'h24;
Memory[8134] = 8'h24;
Memory[8133] = 8'h24;
Memory[8132] = 8'h0B;
Memory[8139] = 8'h1F;
Memory[8138] = 8'h24;
Memory[8137] = 8'h24;
Memory[8136] = 8'h24;
Memory[8143] = 8'h15;
Memory[8142] = 8'h1B;
Memory[8141] = 8'h16;
Memory[8140] = 8'h16;
Memory[8147] = 8'h24;
Memory[8146] = 8'h0A;
Memory[8145] = 8'h16;
Memory[8144] = 8'h0D;
Memory[8151] = 8'h15;
Memory[8150] = 8'h0E;
Memory[8149] = 8'h0E;
Memory[8148] = 8'h24;
Memory[8155] = 8'h1B;
Memory[8154] = 8'h11;
Memory[8153] = 8'h24;
Memory[8152] = 8'h24;
Memory[8159] = 8'h24;
Memory[8158] = 8'h0D;
Memory[8157] = 8'h12;
Memory[8156] = 8'h10;
Memory[8163] = 8'h12;
Memory[8162] = 8'h1C;
Memory[8161] = 8'h0A;
Memory[8160] = 8'h15;
Memory[8167] = 8'h24;
Memory[8166] = 8'h1B;
Memory[8165] = 8'h1F;
Memory[8164] = 8'h1B;
Memory[8171] = 8'h1C;
Memory[8170] = 8'h0E;
Memory[8169] = 8'h16;
Memory[8168] = 8'h16;
Memory[8175] = 8'h1B;
Memory[8174] = 8'h0E;
Memory[8173] = 8'h1C;
Memory[8172] = 8'h1C;
Memory[8179] = 8'h12;
Memory[8178] = 8'h16;
Memory[8177] = 8'h10;
Memory[8176] = 8'h1B;
Memory[8183] = 8'h24;
Memory[8182] = 8'h0B;
Memory[8181] = 8'h1A;
Memory[8180] = 8'h12;
Memory[8187] = 8'h10;
Memory[8186] = 8'h11;
Memory[8185] = 8'h1C;
Memory[8184] = 8'h24;
Memory[8191] = 8'h0B;
Memory[8190] = 8'h1A;
Memory[8189] = 8'h12;
Memory[8188] = 8'h10;
Memory[8195] = 8'h1C;
Memory[8194] = 8'h00;
Memory[8193] = 8'h00;
Memory[8192] = 8'h00;
Memory[8199] = 8'h0B;
Memory[8198] = 8'h1A;
Memory[8197] = 8'h24;
Memory[8196] = 8'h1A;
Memory[8203] = 8'h0A;
Memory[8202] = 8'h16;
Memory[8201] = 8'h10;
Memory[8200] = 8'h0E;
Memory[8207] = 8'h15;
Memory[8206] = 8'h17;
Memory[8205] = 8'h1E;
Memory[8204] = 8'h1E;
Memory[8211] = 8'h24;
Memory[8210] = 8'h00;
Memory[8209] = 8'h00;
Memory[8208] = 8'h00;
Memory[8215] = 8'h11;
Memory[8214] = 8'h12;
Memory[8213] = 8'h10;
Memory[8212] = 8'h11;
Memory[8219] = 8'h24;
Memory[8218] = 8'h00;
Memory[8217] = 8'h00;
Memory[8216] = 8'h00;
Memory[8223] = 8'h15;
Memory[8222] = 8'h0E;
Memory[8221] = 8'h0D;
Memory[8220] = 8'h17;
Memory[8227] = 8'h16;
Memory[8226] = 8'h17;
Memory[8225] = 8'h0F;
Memory[8224] = 8'h0F;
Memory[8231] = 8'h15;
Memory[8230] = 8'h0E;
Memory[8229] = 8'h0D;
Memory[8228] = 8'h24;
Memory[8235] = 8'h24;
Memory[8234] = 8'h17;
Memory[8233] = 8'h16;
Memory[8232] = 8'h24;
Memory[8239] = 8'h15;
Memory[8238] = 8'h0E;
Memory[8237] = 8'h0D;
Memory[8236] = 8'h24;
Memory[8243] = 8'h17;
Memory[8242] = 8'h0F;
Memory[8241] = 8'h0F;
Memory[8240] = 8'h24;
Memory[8247] = 8'h21;
Memory[8246] = 8'h24;
Memory[8245] = 8'h0C;
Memory[8244] = 8'h0A;
Memory[8251] = 8'h16;
Memory[8250] = 8'h17;
Memory[8249] = 8'h16;
Memory[8248] = 8'h24;
Memory[8255] = 8'h24;
Memory[8254] = 8'h0B;
Memory[8253] = 8'h1D;
Memory[8252] = 8'h1B;
Memory[8259] = 8'h14;
Memory[8258] = 8'h0E;
Memory[8257] = 8'h1A;
Memory[8256] = 8'h24;
Memory[8263] = 8'h15;
Memory[8262] = 8'h24;
Memory[8261] = 8'h0E;
Memory[8260] = 8'h0A;
Memory[8267] = 8'h1B;
Memory[8266] = 8'h1F;
Memory[8265] = 8'h24;
Memory[8264] = 8'h15;
Memory[8271] = 8'h21;
Memory[8270] = 8'h24;
Memory[8269] = 8'h11;
Memory[8268] = 8'h0A;
Memory[8275] = 8'h1A;
Memory[8274] = 8'h0D;
Memory[8273] = 8'h24;
Memory[8272] = 8'h21;
Memory[8279] = 8'h22;
Memory[8278] = 8'h22;
Memory[8277] = 8'h22;
Memory[8276] = 8'h22;
Memory[8283] = 8'h22;
Memory[8282] = 8'h22;
Memory[8281] = 8'h01;
Memory[8280] = 8'h22;
Memory[8287] = 8'h22;
Memory[8286] = 8'h22;
Memory[8285] = 8'h22;
Memory[8284] = 8'h22;
Memory[8291] = 8'h01;
Memory[8290] = 8'h22;
Memory[8289] = 8'h08;
Memory[8288] = 8'h08;
Memory[8295] = 8'h24;
Memory[8294] = 8'h24;
Memory[8293] = 8'h18;
Memory[8292] = 8'h0A;
Memory[8299] = 8'h1D;
Memory[8298] = 8'h1B;
Memory[8297] = 8'h0E;
Memory[8296] = 8'h24;
Memory[8303] = 8'h24;
Memory[8302] = 8'h1A;
Memory[8301] = 8'h0E;
Memory[8300] = 8'h1B;
Memory[8307] = 8'h1C;
Memory[8306] = 8'h0A;
Memory[8305] = 8'h1A;
Memory[8304] = 8'h1C;
Memory[8311] = 8'h24;
Memory[8310] = 8'h1A;
Memory[8309] = 8'h0E;
Memory[8308] = 8'h1B;
Memory[8315] = 8'h1D;
Memory[8314] = 8'h16;
Memory[8313] = 8'h16;
Memory[8312] = 8'h0E;
Memory[8319] = 8'h24;
Memory[8318] = 8'h24;
Memory[8317] = 8'h19;
Memory[8316] = 8'h1D;
Memory[8323] = 8'h12;
Memory[8322] = 8'h1C;
Memory[8321] = 8'h24;
Memory[8320] = 8'h24;
Memory[8327] = 8'h16;
Memory[8326] = 8'h16;
Memory[8325] = 8'h1F;
Memory[8324] = 8'h1B;
Memory[8331] = 8'h0C;
Memory[8330] = 8'h17;
Memory[8329] = 8'h1A;
Memory[8328] = 8'h0E;
Memory[8335] = 8'h0C;
Memory[8334] = 8'h17;
Memory[8333] = 8'h16;
Memory[8332] = 8'h10;
Memory[8339] = 8'h1A;
Memory[8338] = 8'h0A;
Memory[8337] = 8'h1C;
Memory[8336] = 8'h0E;
Memory[8343] = 8'h24;
Memory[8342] = 8'h0C;
Memory[8341] = 8'h15;
Memory[8340] = 8'h0E;
Memory[8347] = 8'h0A;
Memory[8346] = 8'h1A;
Memory[8345] = 8'h0E;
Memory[8344] = 8'h0D;
Memory[8351] = 8'h18;
Memory[8350] = 8'h1A;
Memory[8349] = 8'h0E;
Memory[8348] = 8'h1B;
Memory[8355] = 8'h1B;
Memory[8354] = 8'h0A;
Memory[8353] = 8'h16;
Memory[8352] = 8'h1F;
Memory[8359] = 8'h10;
Memory[8358] = 8'h0A;
Memory[8357] = 8'h16;
Memory[8356] = 8'h0E;
Memory[8363] = 8'h17;
Memory[8362] = 8'h1E;
Memory[8361] = 8'h0E;
Memory[8360] = 8'h1A;
Memory[8367] = 8'h24;
Memory[8366] = 8'h24;
Memory[8365] = 8'h00;
Memory[8364] = 8'h00;
Memory[8371] = 8'h00;
Memory[8370] = 8'h00;
Memory[8369] = 8'h00;
Memory[8368] = 8'h00;
Memory[8375] = 8'h1A;
Memory[8374] = 8'h0E;
Memory[8373] = 8'h1B;
Memory[8372] = 8'h0E;
Memory[8379] = 8'h1C;
Memory[8378] = 8'h24;
Memory[8377] = 8'h21;
Memory[8376] = 8'h21;
Memory[8383] = 8'h1A;
Memory[8382] = 8'h0E;
Memory[8381] = 8'h24;
Memory[8380] = 8'h11;
Memory[8387] = 8'h0E;
Memory[8386] = 8'h15;
Memory[8385] = 8'h15;
Memory[8384] = 8'h17;
Memory[8391] = 8'h0A;
Memory[8390] = 8'h16;
Memory[8389] = 8'h18;
Memory[8388] = 8'h15;
Memory[8395] = 8'h1C;
Memory[8394] = 8'h00;
Memory[8393] = 8'h00;
Memory[8392] = 8'h00;
Memory[8399] = 8'h00;
Memory[8398] = 8'h00;
Memory[8397] = 8'h00;
Memory[8396] = 8'h00;
Memory[8403] = 8'h03;
Memory[8402] = 8'h80;
Memory[8401] = 8'h01;
Memory[8400] = 8'h13;
Memory[8407] = 8'h24;
Memory[8406] = 8'h8B;
Memory[8405] = 8'h21;
Memory[8404] = 8'h83;
Memory[8411] = 8'h24;
Memory[8410] = 8'hCB;
Memory[8409] = 8'h22;
Memory[8408] = 8'h03;
Memory[8415] = 8'h01;
Memory[8414] = 8'hA0;
Memory[8413] = 8'h02;
Memory[8412] = 8'h93;
Memory[8419] = 8'h00;
Memory[8418] = 8'h3B;
Memory[8417] = 8'h20;
Memory[8416] = 8'h23;
Memory[8423] = 8'h00;
Memory[8422] = 8'h4B;
Memory[8421] = 8'h22;
Memory[8420] = 8'h23;
Memory[8427] = 8'h00;
Memory[8426] = 8'h5B;
Memory[8425] = 8'h24;
Memory[8424] = 8'h23;
Memory[8431] = 8'h01;
Memory[8430] = 8'hDE;
Memory[8429] = 8'h14;
Memory[8428] = 8'h63;
Memory[8435] = 8'h09;
Memory[8434] = 8'hC0;
Memory[8433] = 8'h00;
Memory[8432] = 8'h6F;
Memory[8439] = 8'h01;
Memory[8438] = 8'hDE;
Memory[8437] = 8'h42;
Memory[8436] = 8'h33;
Memory[8443] = 8'hFF;
Memory[8442] = 8'hF0;
Memory[8441] = 8'h01;
Memory[8440] = 8'h93;
Memory[8447] = 8'h01;
Memory[8446] = 8'hD1;
Memory[8445] = 8'hC1;
Memory[8444] = 8'hB3;
Memory[8451] = 8'h01;
Memory[8450] = 8'h82;
Memory[8449] = 8'h72;
Memory[8448] = 8'h33;
Memory[8455] = 8'h00;
Memory[8454] = 8'h41;
Memory[8453] = 8'hF1;
Memory[8452] = 8'hB3;
Memory[8459] = 8'h00;
Memory[8458] = 8'h01;
Memory[8457] = 8'h94;
Memory[8456] = 8'h63;
Memory[8463] = 8'h2C;
Memory[8462] = 8'h40;
Memory[8461] = 8'h00;
Memory[8460] = 8'h6F;
Memory[8467] = 8'h00;
Memory[8466] = 8'h00;
Memory[8465] = 8'h01;
Memory[8464] = 8'h13;
Memory[8471] = 8'h00;
Memory[8470] = 8'h0E;
Memory[8469] = 8'h8E;
Memory[8468] = 8'h13;
Memory[8475] = 8'h00;
Memory[8474] = 8'h00;
Memory[8473] = 8'h00;
Memory[8472] = 8'h6F;
Memory[8479] = 8'h02;
Memory[8478] = 8'hB0;
Memory[8477] = 8'h01;
Memory[8476] = 8'h93;
Memory[8483] = 8'h00;
Memory[8482] = 8'h31;
Memory[8481] = 8'h06;
Memory[8480] = 8'h63;
Memory[8487] = 8'h00;
Memory[8486] = 8'h0F;
Memory[8485] = 8'h8F;
Memory[8484] = 8'h13;
Memory[8491] = 8'h09;
Memory[8490] = 8'hC0;
Memory[8489] = 8'h00;
Memory[8488] = 8'h6F;
Memory[8495] = 8'h26;
Memory[8494] = 8'h0B;
Memory[8493] = 8'h21;
Memory[8492] = 8'h83;
Memory[8499] = 8'h00;
Memory[8498] = 8'h10;
Memory[8497] = 8'h02;
Memory[8496] = 8'h13;
Memory[8503] = 8'h00;
Memory[8502] = 8'h41;
Memory[8501] = 8'h84;
Memory[8500] = 8'h63;
Memory[8507] = 8'h12;
Memory[8506] = 8'h40;
Memory[8505] = 8'h20;
Memory[8504] = 8'h6F;
Memory[8511] = 8'h05;
Memory[8510] = 8'h0B;
Memory[8509] = 8'h22;
Memory[8508] = 8'h03;
Memory[8515] = 8'h40;
Memory[8514] = 8'h4F;
Memory[8513] = 8'h81;
Memory[8512] = 8'hB3;
Memory[8519] = 8'h05;
Memory[8518] = 8'h4B;
Memory[8517] = 8'h22;
Memory[8516] = 8'h03;
Memory[8523] = 8'h00;
Memory[8522] = 8'h32;
Memory[8521] = 8'h22;
Memory[8520] = 8'hB3;
Memory[8527] = 8'h00;
Memory[8526] = 8'h02;
Memory[8525] = 8'h84;
Memory[8524] = 8'h63;
Memory[8531] = 8'h78;
Memory[8530] = 8'h10;
Memory[8529] = 8'h50;
Memory[8528] = 8'h6F;
Memory[8535] = 8'h6E;
Memory[8534] = 8'h4C;
Memory[8533] = 8'hA2;
Memory[8532] = 8'h03;
Memory[8539] = 8'h00;
Memory[8538] = 8'h32;
Memory[8537] = 8'h22;
Memory[8536] = 8'hB3;
Memory[8543] = 8'h00;
Memory[8542] = 8'h02;
Memory[8541] = 8'h84;
Memory[8540] = 8'h63;
Memory[8547] = 8'h77;
Memory[8546] = 8'h50;
Memory[8545] = 8'h50;
Memory[8544] = 8'h6F;
Memory[8551] = 8'h6E;
Memory[8550] = 8'h0C;
Memory[8549] = 8'hA2;
Memory[8548] = 8'h03;
Memory[8555] = 8'h00;
Memory[8554] = 8'h32;
Memory[8553] = 8'h22;
Memory[8552] = 8'hB3;
Memory[8559] = 8'h00;
Memory[8558] = 8'h02;
Memory[8557] = 8'h84;
Memory[8556] = 8'h63;
Memory[8563] = 8'h76;
Memory[8562] = 8'h90;
Memory[8561] = 8'h50;
Memory[8560] = 8'h6F;
Memory[8567] = 8'h6D;
Memory[8566] = 8'hCC;
Memory[8565] = 8'hA2;
Memory[8564] = 8'h03;
Memory[8571] = 8'h00;
Memory[8570] = 8'h32;
Memory[8569] = 8'h22;
Memory[8568] = 8'hB3;
Memory[8575] = 8'h00;
Memory[8574] = 8'h02;
Memory[8573] = 8'h84;
Memory[8572] = 8'h63;
Memory[8579] = 8'h75;
Memory[8578] = 8'hD0;
Memory[8577] = 8'h50;
Memory[8576] = 8'h6F;
Memory[8583] = 8'h6D;
Memory[8582] = 8'h8C;
Memory[8581] = 8'hA2;
Memory[8580] = 8'h03;
Memory[8587] = 8'h00;
Memory[8586] = 8'h32;
Memory[8585] = 8'h22;
Memory[8584] = 8'hB3;
Memory[8591] = 8'h00;
Memory[8590] = 8'h02;
Memory[8589] = 8'h84;
Memory[8588] = 8'h63;
Memory[8595] = 8'h75;
Memory[8594] = 8'h10;
Memory[8593] = 8'h50;
Memory[8592] = 8'h6F;
Memory[8599] = 8'h6D;
Memory[8598] = 8'h4C;
Memory[8597] = 8'hA2;
Memory[8596] = 8'h03;
Memory[8603] = 8'h00;
Memory[8602] = 8'h32;
Memory[8601] = 8'h22;
Memory[8600] = 8'hB3;
Memory[8607] = 8'h00;
Memory[8606] = 8'h02;
Memory[8605] = 8'h84;
Memory[8604] = 8'h63;
Memory[8611] = 8'h74;
Memory[8610] = 8'h50;
Memory[8609] = 8'h50;
Memory[8608] = 8'h6F;
Memory[8615] = 8'h6D;
Memory[8614] = 8'h0C;
Memory[8613] = 8'hA2;
Memory[8612] = 8'h03;
Memory[8619] = 8'h00;
Memory[8618] = 8'h32;
Memory[8617] = 8'h22;
Memory[8616] = 8'hB3;
Memory[8623] = 8'h00;
Memory[8622] = 8'h02;
Memory[8621] = 8'h84;
Memory[8620] = 8'h63;
Memory[8627] = 8'h73;
Memory[8626] = 8'h90;
Memory[8625] = 8'h50;
Memory[8624] = 8'h6F;
Memory[8631] = 8'h6C;
Memory[8630] = 8'hCC;
Memory[8629] = 8'hA2;
Memory[8628] = 8'h03;
Memory[8635] = 8'h00;
Memory[8634] = 8'h32;
Memory[8633] = 8'h22;
Memory[8632] = 8'hB3;
Memory[8639] = 8'h00;
Memory[8638] = 8'h02;
Memory[8637] = 8'h84;
Memory[8636] = 8'h63;
Memory[8643] = 8'h72;
Memory[8642] = 8'hD0;
Memory[8641] = 8'h50;
Memory[8640] = 8'h6F;
Memory[8647] = 8'h6C;
Memory[8646] = 8'h8C;
Memory[8645] = 8'hA2;
Memory[8644] = 8'h03;
Memory[8651] = 8'h00;
Memory[8650] = 8'h32;
Memory[8649] = 8'h22;
Memory[8648] = 8'hB3;
Memory[8655] = 8'h00;
Memory[8654] = 8'h02;
Memory[8653] = 8'h84;
Memory[8652] = 8'h63;
Memory[8659] = 8'h72;
Memory[8658] = 8'h10;
Memory[8657] = 8'h50;
Memory[8656] = 8'h6F;
Memory[8663] = 8'h6C;
Memory[8662] = 8'h4C;
Memory[8661] = 8'hA2;
Memory[8660] = 8'h03;
Memory[8667] = 8'h00;
Memory[8666] = 8'h32;
Memory[8665] = 8'h22;
Memory[8664] = 8'hB3;
Memory[8671] = 8'h00;
Memory[8670] = 8'h02;
Memory[8669] = 8'h84;
Memory[8668] = 8'h63;
Memory[8675] = 8'h71;
Memory[8674] = 8'h50;
Memory[8673] = 8'h50;
Memory[8672] = 8'h6F;
Memory[8679] = 8'h6C;
Memory[8678] = 8'h0C;
Memory[8677] = 8'hA2;
Memory[8676] = 8'h03;
Memory[8683] = 8'h00;
Memory[8682] = 8'h32;
Memory[8681] = 8'h22;
Memory[8680] = 8'hB3;
Memory[8687] = 8'h00;
Memory[8686] = 8'h02;
Memory[8685] = 8'h84;
Memory[8684] = 8'h63;
Memory[8691] = 8'h70;
Memory[8690] = 8'h90;
Memory[8689] = 8'h50;
Memory[8688] = 8'h6F;
Memory[8695] = 8'h6B;
Memory[8694] = 8'hCC;
Memory[8693] = 8'hA2;
Memory[8692] = 8'h03;
Memory[8699] = 8'h00;
Memory[8698] = 8'h32;
Memory[8697] = 8'h22;
Memory[8696] = 8'hB3;
Memory[8703] = 8'h00;
Memory[8702] = 8'h02;
Memory[8701] = 8'h84;
Memory[8700] = 8'h63;
Memory[8707] = 8'h6F;
Memory[8706] = 8'hD0;
Memory[8705] = 8'h50;
Memory[8704] = 8'h6F;
Memory[8711] = 8'h6B;
Memory[8710] = 8'h8C;
Memory[8709] = 8'hA2;
Memory[8708] = 8'h03;
Memory[8715] = 8'h00;
Memory[8714] = 8'h32;
Memory[8713] = 8'h22;
Memory[8712] = 8'hB3;
Memory[8719] = 8'h00;
Memory[8718] = 8'h02;
Memory[8717] = 8'h84;
Memory[8716] = 8'h63;
Memory[8723] = 8'h6F;
Memory[8722] = 8'h10;
Memory[8721] = 8'h50;
Memory[8720] = 8'h6F;
Memory[8727] = 8'h6B;
Memory[8726] = 8'h4C;
Memory[8725] = 8'hA2;
Memory[8724] = 8'h03;
Memory[8731] = 8'h00;
Memory[8730] = 8'h32;
Memory[8729] = 8'h22;
Memory[8728] = 8'hB3;
Memory[8735] = 8'h00;
Memory[8734] = 8'h02;
Memory[8733] = 8'h84;
Memory[8732] = 8'h63;
Memory[8739] = 8'h6E;
Memory[8738] = 8'h50;
Memory[8737] = 8'h50;
Memory[8736] = 8'h6F;
Memory[8743] = 8'h6B;
Memory[8742] = 8'h0C;
Memory[8741] = 8'hA2;
Memory[8740] = 8'h03;
Memory[8747] = 8'h00;
Memory[8746] = 8'h32;
Memory[8745] = 8'h22;
Memory[8744] = 8'hB3;
Memory[8751] = 8'h00;
Memory[8750] = 8'h02;
Memory[8749] = 8'h84;
Memory[8748] = 8'h63;
Memory[8755] = 8'h6D;
Memory[8754] = 8'h90;
Memory[8753] = 8'h50;
Memory[8752] = 8'h6F;
Memory[8759] = 8'h6A;
Memory[8758] = 8'hCC;
Memory[8757] = 8'hA2;
Memory[8756] = 8'h03;
Memory[8763] = 8'h00;
Memory[8762] = 8'h32;
Memory[8761] = 8'h22;
Memory[8760] = 8'hB3;
Memory[8767] = 8'h00;
Memory[8766] = 8'h02;
Memory[8765] = 8'h84;
Memory[8764] = 8'h63;
Memory[8771] = 8'h6C;
Memory[8770] = 8'hD0;
Memory[8769] = 8'h50;
Memory[8768] = 8'h6F;
Memory[8775] = 8'h6A;
Memory[8774] = 8'h8C;
Memory[8773] = 8'hA2;
Memory[8772] = 8'h03;
Memory[8779] = 8'h00;
Memory[8778] = 8'h32;
Memory[8777] = 8'h22;
Memory[8776] = 8'hB3;
Memory[8783] = 8'h00;
Memory[8782] = 8'h02;
Memory[8781] = 8'h84;
Memory[8780] = 8'h63;
Memory[8787] = 8'h6C;
Memory[8786] = 8'h10;
Memory[8785] = 8'h50;
Memory[8784] = 8'h6F;
Memory[8791] = 8'h6A;
Memory[8790] = 8'h4C;
Memory[8789] = 8'hA2;
Memory[8788] = 8'h03;
Memory[8795] = 8'h00;
Memory[8794] = 8'h32;
Memory[8793] = 8'h22;
Memory[8792] = 8'hB3;
Memory[8799] = 8'h00;
Memory[8798] = 8'h02;
Memory[8797] = 8'h84;
Memory[8796] = 8'h63;
Memory[8803] = 8'h6B;
Memory[8802] = 8'h50;
Memory[8801] = 8'h50;
Memory[8800] = 8'h6F;
Memory[8807] = 8'h6A;
Memory[8806] = 8'h0C;
Memory[8805] = 8'hA2;
Memory[8804] = 8'h03;
Memory[8811] = 8'h00;
Memory[8810] = 8'h32;
Memory[8809] = 8'h22;
Memory[8808] = 8'hB3;
Memory[8815] = 8'h00;
Memory[8814] = 8'h02;
Memory[8813] = 8'h84;
Memory[8812] = 8'h63;
Memory[8819] = 8'h6A;
Memory[8818] = 8'h90;
Memory[8817] = 8'h50;
Memory[8816] = 8'h6F;
Memory[8823] = 8'h69;
Memory[8822] = 8'hCC;
Memory[8821] = 8'hA2;
Memory[8820] = 8'h03;
Memory[8827] = 8'h00;
Memory[8826] = 8'h32;
Memory[8825] = 8'h22;
Memory[8824] = 8'hB3;
Memory[8831] = 8'h00;
Memory[8830] = 8'h02;
Memory[8829] = 8'h84;
Memory[8828] = 8'h63;
Memory[8835] = 8'h69;
Memory[8834] = 8'hD0;
Memory[8833] = 8'h50;
Memory[8832] = 8'h6F;
Memory[8839] = 8'h69;
Memory[8838] = 8'h8C;
Memory[8837] = 8'hA2;
Memory[8836] = 8'h03;
Memory[8843] = 8'h00;
Memory[8842] = 8'h32;
Memory[8841] = 8'h22;
Memory[8840] = 8'hB3;
Memory[8847] = 8'h00;
Memory[8846] = 8'h02;
Memory[8845] = 8'h84;
Memory[8844] = 8'h63;
Memory[8851] = 8'h69;
Memory[8850] = 8'h10;
Memory[8849] = 8'h50;
Memory[8848] = 8'h6F;
Memory[8855] = 8'h69;
Memory[8854] = 8'h4C;
Memory[8853] = 8'hA2;
Memory[8852] = 8'h03;
Memory[8859] = 8'h00;
Memory[8858] = 8'h32;
Memory[8857] = 8'h22;
Memory[8856] = 8'hB3;
Memory[8863] = 8'h00;
Memory[8862] = 8'h02;
Memory[8861] = 8'h84;
Memory[8860] = 8'h63;
Memory[8867] = 8'h68;
Memory[8866] = 8'h50;
Memory[8865] = 8'h50;
Memory[8864] = 8'h6F;
Memory[8871] = 8'h69;
Memory[8870] = 8'h0C;
Memory[8869] = 8'hA2;
Memory[8868] = 8'h03;
Memory[8875] = 8'h00;
Memory[8874] = 8'h32;
Memory[8873] = 8'h22;
Memory[8872] = 8'hB3;
Memory[8879] = 8'h00;
Memory[8878] = 8'h02;
Memory[8877] = 8'h84;
Memory[8876] = 8'h63;
Memory[8883] = 8'h67;
Memory[8882] = 8'h90;
Memory[8881] = 8'h50;
Memory[8880] = 8'h6F;
Memory[8887] = 8'h68;
Memory[8886] = 8'hCC;
Memory[8885] = 8'hA2;
Memory[8884] = 8'h03;
Memory[8891] = 8'h00;
Memory[8890] = 8'h32;
Memory[8889] = 8'h22;
Memory[8888] = 8'hB3;
Memory[8895] = 8'h00;
Memory[8894] = 8'h02;
Memory[8893] = 8'h84;
Memory[8892] = 8'h63;
Memory[8899] = 8'h66;
Memory[8898] = 8'hD0;
Memory[8897] = 8'h50;
Memory[8896] = 8'h6F;
Memory[8903] = 8'h68;
Memory[8902] = 8'h8C;
Memory[8901] = 8'hA2;
Memory[8900] = 8'h03;
Memory[8907] = 8'h00;
Memory[8906] = 8'h32;
Memory[8905] = 8'h22;
Memory[8904] = 8'hB3;
Memory[8911] = 8'h00;
Memory[8910] = 8'h02;
Memory[8909] = 8'h84;
Memory[8908] = 8'h63;
Memory[8915] = 8'h66;
Memory[8914] = 8'h10;
Memory[8913] = 8'h50;
Memory[8912] = 8'h6F;
Memory[8919] = 8'h68;
Memory[8918] = 8'h4C;
Memory[8917] = 8'hA2;
Memory[8916] = 8'h03;
Memory[8923] = 8'h00;
Memory[8922] = 8'h32;
Memory[8921] = 8'h22;
Memory[8920] = 8'hB3;
Memory[8927] = 8'h00;
Memory[8926] = 8'h02;
Memory[8925] = 8'h84;
Memory[8924] = 8'h63;
Memory[8931] = 8'h65;
Memory[8930] = 8'h50;
Memory[8929] = 8'h50;
Memory[8928] = 8'h6F;
Memory[8935] = 8'h68;
Memory[8934] = 8'h0C;
Memory[8933] = 8'hA2;
Memory[8932] = 8'h03;
Memory[8939] = 8'h00;
Memory[8938] = 8'h32;
Memory[8937] = 8'h22;
Memory[8936] = 8'hB3;
Memory[8943] = 8'h00;
Memory[8942] = 8'h02;
Memory[8941] = 8'h84;
Memory[8940] = 8'h63;
Memory[8947] = 8'h64;
Memory[8946] = 8'h90;
Memory[8945] = 8'h50;
Memory[8944] = 8'h6F;
Memory[8951] = 8'h67;
Memory[8950] = 8'hCC;
Memory[8949] = 8'hA2;
Memory[8948] = 8'h03;
Memory[8955] = 8'h00;
Memory[8954] = 8'h32;
Memory[8953] = 8'h22;
Memory[8952] = 8'hB3;
Memory[8959] = 8'h00;
Memory[8958] = 8'h02;
Memory[8957] = 8'h84;
Memory[8956] = 8'h63;
Memory[8963] = 8'h63;
Memory[8962] = 8'hD0;
Memory[8961] = 8'h50;
Memory[8960] = 8'h6F;
Memory[8967] = 8'h67;
Memory[8966] = 8'h8C;
Memory[8965] = 8'hA2;
Memory[8964] = 8'h03;
Memory[8971] = 8'h00;
Memory[8970] = 8'h32;
Memory[8969] = 8'h22;
Memory[8968] = 8'hB3;
Memory[8975] = 8'h00;
Memory[8974] = 8'h02;
Memory[8973] = 8'h84;
Memory[8972] = 8'h63;
Memory[8979] = 8'h63;
Memory[8978] = 8'h10;
Memory[8977] = 8'h50;
Memory[8976] = 8'h6F;
Memory[8983] = 8'h67;
Memory[8982] = 8'h4C;
Memory[8981] = 8'hA2;
Memory[8980] = 8'h03;
Memory[8987] = 8'h00;
Memory[8986] = 8'h32;
Memory[8985] = 8'h22;
Memory[8984] = 8'hB3;
Memory[8991] = 8'h00;
Memory[8990] = 8'h02;
Memory[8989] = 8'h84;
Memory[8988] = 8'h63;
Memory[8995] = 8'h62;
Memory[8994] = 8'h50;
Memory[8993] = 8'h50;
Memory[8992] = 8'h6F;
Memory[8999] = 8'h67;
Memory[8998] = 8'h0C;
Memory[8997] = 8'hA2;
Memory[8996] = 8'h03;
Memory[9003] = 8'h00;
Memory[9002] = 8'h32;
Memory[9001] = 8'h22;
Memory[9000] = 8'hB3;
Memory[9007] = 8'h00;
Memory[9006] = 8'h02;
Memory[9005] = 8'h84;
Memory[9004] = 8'h63;
Memory[9011] = 8'h61;
Memory[9010] = 8'h90;
Memory[9009] = 8'h50;
Memory[9008] = 8'h6F;
Memory[9015] = 8'h66;
Memory[9014] = 8'hCC;
Memory[9013] = 8'hA2;
Memory[9012] = 8'h03;
Memory[9019] = 8'h00;
Memory[9018] = 8'h32;
Memory[9017] = 8'h22;
Memory[9016] = 8'hB3;
Memory[9023] = 8'h00;
Memory[9022] = 8'h02;
Memory[9021] = 8'h84;
Memory[9020] = 8'h63;
Memory[9027] = 8'h60;
Memory[9026] = 8'hD0;
Memory[9025] = 8'h50;
Memory[9024] = 8'h6F;
Memory[9031] = 8'h66;
Memory[9030] = 8'h8C;
Memory[9029] = 8'hA2;
Memory[9028] = 8'h03;
Memory[9035] = 8'h00;
Memory[9034] = 8'h32;
Memory[9033] = 8'h22;
Memory[9032] = 8'hB3;
Memory[9039] = 8'h00;
Memory[9038] = 8'h02;
Memory[9037] = 8'h84;
Memory[9036] = 8'h63;
Memory[9043] = 8'h60;
Memory[9042] = 8'h10;
Memory[9041] = 8'h50;
Memory[9040] = 8'h6F;
Memory[9047] = 8'h66;
Memory[9046] = 8'h4C;
Memory[9045] = 8'hA2;
Memory[9044] = 8'h03;
Memory[9051] = 8'h00;
Memory[9050] = 8'h32;
Memory[9049] = 8'h22;
Memory[9048] = 8'hB3;
Memory[9055] = 8'h00;
Memory[9054] = 8'h02;
Memory[9053] = 8'h84;
Memory[9052] = 8'h63;
Memory[9059] = 8'h5F;
Memory[9058] = 8'h50;
Memory[9057] = 8'h50;
Memory[9056] = 8'h6F;
Memory[9063] = 8'h66;
Memory[9062] = 8'h0C;
Memory[9061] = 8'hA2;
Memory[9060] = 8'h03;
Memory[9067] = 8'h00;
Memory[9066] = 8'h32;
Memory[9065] = 8'h22;
Memory[9064] = 8'hB3;
Memory[9071] = 8'h00;
Memory[9070] = 8'h02;
Memory[9069] = 8'h84;
Memory[9068] = 8'h63;
Memory[9075] = 8'h5E;
Memory[9074] = 8'h90;
Memory[9073] = 8'h50;
Memory[9072] = 8'h6F;
Memory[9079] = 8'h65;
Memory[9078] = 8'hCC;
Memory[9077] = 8'hA2;
Memory[9076] = 8'h03;
Memory[9083] = 8'h00;
Memory[9082] = 8'h32;
Memory[9081] = 8'h22;
Memory[9080] = 8'hB3;
Memory[9087] = 8'h00;
Memory[9086] = 8'h02;
Memory[9085] = 8'h84;
Memory[9084] = 8'h63;
Memory[9091] = 8'h5D;
Memory[9090] = 8'hD0;
Memory[9089] = 8'h50;
Memory[9088] = 8'h6F;
Memory[9095] = 8'h65;
Memory[9094] = 8'h8C;
Memory[9093] = 8'hA2;
Memory[9092] = 8'h03;
Memory[9099] = 8'h00;
Memory[9098] = 8'h32;
Memory[9097] = 8'h22;
Memory[9096] = 8'hB3;
Memory[9103] = 8'h00;
Memory[9102] = 8'h02;
Memory[9101] = 8'h84;
Memory[9100] = 8'h63;
Memory[9107] = 8'h5D;
Memory[9106] = 8'h10;
Memory[9105] = 8'h50;
Memory[9104] = 8'h6F;
Memory[9111] = 8'h65;
Memory[9110] = 8'h4C;
Memory[9109] = 8'hA2;
Memory[9108] = 8'h03;
Memory[9115] = 8'h00;
Memory[9114] = 8'h32;
Memory[9113] = 8'h22;
Memory[9112] = 8'hB3;
Memory[9119] = 8'h00;
Memory[9118] = 8'h02;
Memory[9117] = 8'h84;
Memory[9116] = 8'h63;
Memory[9123] = 8'h5C;
Memory[9122] = 8'h50;
Memory[9121] = 8'h50;
Memory[9120] = 8'h6F;
Memory[9127] = 8'h65;
Memory[9126] = 8'h0C;
Memory[9125] = 8'hA2;
Memory[9124] = 8'h03;
Memory[9131] = 8'h00;
Memory[9130] = 8'h32;
Memory[9129] = 8'h22;
Memory[9128] = 8'hB3;
Memory[9135] = 8'h00;
Memory[9134] = 8'h02;
Memory[9133] = 8'h84;
Memory[9132] = 8'h63;
Memory[9139] = 8'h5B;
Memory[9138] = 8'h90;
Memory[9137] = 8'h50;
Memory[9136] = 8'h6F;
Memory[9143] = 8'h64;
Memory[9142] = 8'hCC;
Memory[9141] = 8'hA2;
Memory[9140] = 8'h03;
Memory[9147] = 8'h00;
Memory[9146] = 8'h32;
Memory[9145] = 8'h22;
Memory[9144] = 8'hB3;
Memory[9151] = 8'h00;
Memory[9150] = 8'h02;
Memory[9149] = 8'h84;
Memory[9148] = 8'h63;
Memory[9155] = 8'h5A;
Memory[9154] = 8'hD0;
Memory[9153] = 8'h50;
Memory[9152] = 8'h6F;
Memory[9159] = 8'h64;
Memory[9158] = 8'h8C;
Memory[9157] = 8'hA2;
Memory[9156] = 8'h03;
Memory[9163] = 8'h00;
Memory[9162] = 8'h32;
Memory[9161] = 8'h22;
Memory[9160] = 8'hB3;
Memory[9167] = 8'h00;
Memory[9166] = 8'h02;
Memory[9165] = 8'h84;
Memory[9164] = 8'h63;
Memory[9171] = 8'h5A;
Memory[9170] = 8'h10;
Memory[9169] = 8'h50;
Memory[9168] = 8'h6F;
Memory[9175] = 8'h64;
Memory[9174] = 8'h4C;
Memory[9173] = 8'hA2;
Memory[9172] = 8'h03;
Memory[9179] = 8'h00;
Memory[9178] = 8'h32;
Memory[9177] = 8'h22;
Memory[9176] = 8'hB3;
Memory[9183] = 8'h00;
Memory[9182] = 8'h02;
Memory[9181] = 8'h84;
Memory[9180] = 8'h63;
Memory[9187] = 8'h59;
Memory[9186] = 8'h50;
Memory[9185] = 8'h50;
Memory[9184] = 8'h6F;
Memory[9191] = 8'h64;
Memory[9190] = 8'h0C;
Memory[9189] = 8'hA2;
Memory[9188] = 8'h03;
Memory[9195] = 8'h00;
Memory[9194] = 8'h32;
Memory[9193] = 8'h22;
Memory[9192] = 8'hB3;
Memory[9199] = 8'h00;
Memory[9198] = 8'h02;
Memory[9197] = 8'h84;
Memory[9196] = 8'h63;
Memory[9203] = 8'h58;
Memory[9202] = 8'h90;
Memory[9201] = 8'h50;
Memory[9200] = 8'h6F;
Memory[9207] = 8'h63;
Memory[9206] = 8'hCC;
Memory[9205] = 8'hA2;
Memory[9204] = 8'h03;
Memory[9211] = 8'h00;
Memory[9210] = 8'h32;
Memory[9209] = 8'h22;
Memory[9208] = 8'hB3;
Memory[9215] = 8'h00;
Memory[9214] = 8'h02;
Memory[9213] = 8'h84;
Memory[9212] = 8'h63;
Memory[9219] = 8'h57;
Memory[9218] = 8'hD0;
Memory[9217] = 8'h50;
Memory[9216] = 8'h6F;
Memory[9223] = 8'h63;
Memory[9222] = 8'h8C;
Memory[9221] = 8'hA2;
Memory[9220] = 8'h03;
Memory[9227] = 8'h00;
Memory[9226] = 8'h32;
Memory[9225] = 8'h22;
Memory[9224] = 8'hB3;
Memory[9231] = 8'h00;
Memory[9230] = 8'h02;
Memory[9229] = 8'h84;
Memory[9228] = 8'h63;
Memory[9235] = 8'h57;
Memory[9234] = 8'h10;
Memory[9233] = 8'h50;
Memory[9232] = 8'h6F;
Memory[9239] = 8'h63;
Memory[9238] = 8'h4C;
Memory[9237] = 8'hA2;
Memory[9236] = 8'h03;
Memory[9243] = 8'h00;
Memory[9242] = 8'h32;
Memory[9241] = 8'h22;
Memory[9240] = 8'hB3;
Memory[9247] = 8'h00;
Memory[9246] = 8'h02;
Memory[9245] = 8'h84;
Memory[9244] = 8'h63;
Memory[9251] = 8'h56;
Memory[9250] = 8'h50;
Memory[9249] = 8'h50;
Memory[9248] = 8'h6F;
Memory[9255] = 8'h63;
Memory[9254] = 8'h0C;
Memory[9253] = 8'hA2;
Memory[9252] = 8'h03;
Memory[9259] = 8'h00;
Memory[9258] = 8'h32;
Memory[9257] = 8'h22;
Memory[9256] = 8'hB3;
Memory[9263] = 8'h00;
Memory[9262] = 8'h02;
Memory[9261] = 8'h84;
Memory[9260] = 8'h63;
Memory[9267] = 8'h55;
Memory[9266] = 8'h90;
Memory[9265] = 8'h50;
Memory[9264] = 8'h6F;
Memory[9271] = 8'h62;
Memory[9270] = 8'hCC;
Memory[9269] = 8'hA2;
Memory[9268] = 8'h03;
Memory[9275] = 8'h00;
Memory[9274] = 8'h32;
Memory[9273] = 8'h22;
Memory[9272] = 8'hB3;
Memory[9279] = 8'h00;
Memory[9278] = 8'h02;
Memory[9277] = 8'h84;
Memory[9276] = 8'h63;
Memory[9283] = 8'h54;
Memory[9282] = 8'hD0;
Memory[9281] = 8'h50;
Memory[9280] = 8'h6F;
Memory[9287] = 8'h62;
Memory[9286] = 8'h8C;
Memory[9285] = 8'hA2;
Memory[9284] = 8'h03;
Memory[9291] = 8'h00;
Memory[9290] = 8'h32;
Memory[9289] = 8'h22;
Memory[9288] = 8'hB3;
Memory[9295] = 8'h00;
Memory[9294] = 8'h02;
Memory[9293] = 8'h84;
Memory[9292] = 8'h63;
Memory[9299] = 8'h54;
Memory[9298] = 8'h10;
Memory[9297] = 8'h50;
Memory[9296] = 8'h6F;
Memory[9303] = 8'h62;
Memory[9302] = 8'h4C;
Memory[9301] = 8'hA2;
Memory[9300] = 8'h03;
Memory[9307] = 8'h00;
Memory[9306] = 8'h32;
Memory[9305] = 8'h22;
Memory[9304] = 8'hB3;
Memory[9311] = 8'h00;
Memory[9310] = 8'h02;
Memory[9309] = 8'h84;
Memory[9308] = 8'h63;
Memory[9315] = 8'h53;
Memory[9314] = 8'h50;
Memory[9313] = 8'h50;
Memory[9312] = 8'h6F;
Memory[9319] = 8'h62;
Memory[9318] = 8'h0C;
Memory[9317] = 8'hA2;
Memory[9316] = 8'h03;
Memory[9323] = 8'h00;
Memory[9322] = 8'h32;
Memory[9321] = 8'h22;
Memory[9320] = 8'hB3;
Memory[9327] = 8'h00;
Memory[9326] = 8'h02;
Memory[9325] = 8'h84;
Memory[9324] = 8'h63;
Memory[9331] = 8'h52;
Memory[9330] = 8'h90;
Memory[9329] = 8'h50;
Memory[9328] = 8'h6F;
Memory[9335] = 8'h61;
Memory[9334] = 8'hCC;
Memory[9333] = 8'hA2;
Memory[9332] = 8'h03;
Memory[9339] = 8'h00;
Memory[9338] = 8'h32;
Memory[9337] = 8'h22;
Memory[9336] = 8'hB3;
Memory[9343] = 8'h00;
Memory[9342] = 8'h02;
Memory[9341] = 8'h84;
Memory[9340] = 8'h63;
Memory[9347] = 8'h51;
Memory[9346] = 8'hD0;
Memory[9345] = 8'h50;
Memory[9344] = 8'h6F;
Memory[9351] = 8'h61;
Memory[9350] = 8'h8C;
Memory[9349] = 8'hA2;
Memory[9348] = 8'h03;
Memory[9355] = 8'h00;
Memory[9354] = 8'h32;
Memory[9353] = 8'h22;
Memory[9352] = 8'hB3;
Memory[9359] = 8'h00;
Memory[9358] = 8'h02;
Memory[9357] = 8'h84;
Memory[9356] = 8'h63;
Memory[9363] = 8'h51;
Memory[9362] = 8'h10;
Memory[9361] = 8'h50;
Memory[9360] = 8'h6F;
Memory[9367] = 8'h61;
Memory[9366] = 8'h4C;
Memory[9365] = 8'hA2;
Memory[9364] = 8'h03;
Memory[9371] = 8'h00;
Memory[9370] = 8'h32;
Memory[9369] = 8'h22;
Memory[9368] = 8'hB3;
Memory[9375] = 8'h00;
Memory[9374] = 8'h02;
Memory[9373] = 8'h84;
Memory[9372] = 8'h63;
Memory[9379] = 8'h50;
Memory[9378] = 8'h50;
Memory[9377] = 8'h50;
Memory[9376] = 8'h6F;
Memory[9383] = 8'h61;
Memory[9382] = 8'h0C;
Memory[9381] = 8'hA2;
Memory[9380] = 8'h03;
Memory[9387] = 8'h00;
Memory[9386] = 8'h32;
Memory[9385] = 8'h22;
Memory[9384] = 8'hB3;
Memory[9391] = 8'h00;
Memory[9390] = 8'h02;
Memory[9389] = 8'h84;
Memory[9388] = 8'h63;
Memory[9395] = 8'h4F;
Memory[9394] = 8'h90;
Memory[9393] = 8'h50;
Memory[9392] = 8'h6F;
Memory[9399] = 8'h60;
Memory[9398] = 8'hCC;
Memory[9397] = 8'hA2;
Memory[9396] = 8'h03;
Memory[9403] = 8'h00;
Memory[9402] = 8'h32;
Memory[9401] = 8'h22;
Memory[9400] = 8'hB3;
Memory[9407] = 8'h00;
Memory[9406] = 8'h02;
Memory[9405] = 8'h84;
Memory[9404] = 8'h63;
Memory[9411] = 8'h4E;
Memory[9410] = 8'hD0;
Memory[9409] = 8'h50;
Memory[9408] = 8'h6F;
Memory[9415] = 8'h60;
Memory[9414] = 8'h8C;
Memory[9413] = 8'hA2;
Memory[9412] = 8'h03;
Memory[9419] = 8'h00;
Memory[9418] = 8'h32;
Memory[9417] = 8'h22;
Memory[9416] = 8'hB3;
Memory[9423] = 8'h00;
Memory[9422] = 8'h02;
Memory[9421] = 8'h84;
Memory[9420] = 8'h63;
Memory[9427] = 8'h4E;
Memory[9426] = 8'h10;
Memory[9425] = 8'h50;
Memory[9424] = 8'h6F;
Memory[9431] = 8'h60;
Memory[9430] = 8'h4C;
Memory[9429] = 8'hA2;
Memory[9428] = 8'h03;
Memory[9435] = 8'h00;
Memory[9434] = 8'h32;
Memory[9433] = 8'h22;
Memory[9432] = 8'hB3;
Memory[9439] = 8'h00;
Memory[9438] = 8'h02;
Memory[9437] = 8'h84;
Memory[9436] = 8'h63;
Memory[9443] = 8'h4D;
Memory[9442] = 8'h50;
Memory[9441] = 8'h50;
Memory[9440] = 8'h6F;
Memory[9447] = 8'h60;
Memory[9446] = 8'h0C;
Memory[9445] = 8'hA2;
Memory[9444] = 8'h03;
Memory[9451] = 8'h00;
Memory[9450] = 8'h32;
Memory[9449] = 8'h22;
Memory[9448] = 8'hB3;
Memory[9455] = 8'h00;
Memory[9454] = 8'h02;
Memory[9453] = 8'h84;
Memory[9452] = 8'h63;
Memory[9459] = 8'h4C;
Memory[9458] = 8'h90;
Memory[9457] = 8'h50;
Memory[9456] = 8'h6F;
Memory[9463] = 8'h5F;
Memory[9462] = 8'hCC;
Memory[9461] = 8'hA2;
Memory[9460] = 8'h03;
Memory[9467] = 8'h00;
Memory[9466] = 8'h32;
Memory[9465] = 8'h22;
Memory[9464] = 8'hB3;
Memory[9471] = 8'h00;
Memory[9470] = 8'h02;
Memory[9469] = 8'h84;
Memory[9468] = 8'h63;
Memory[9475] = 8'h4B;
Memory[9474] = 8'hD0;
Memory[9473] = 8'h50;
Memory[9472] = 8'h6F;
Memory[9479] = 8'h5F;
Memory[9478] = 8'h8C;
Memory[9477] = 8'hA2;
Memory[9476] = 8'h03;
Memory[9483] = 8'h00;
Memory[9482] = 8'h32;
Memory[9481] = 8'h22;
Memory[9480] = 8'hB3;
Memory[9487] = 8'h00;
Memory[9486] = 8'h02;
Memory[9485] = 8'h84;
Memory[9484] = 8'h63;
Memory[9491] = 8'h4B;
Memory[9490] = 8'h10;
Memory[9489] = 8'h50;
Memory[9488] = 8'h6F;
Memory[9495] = 8'h5F;
Memory[9494] = 8'h4C;
Memory[9493] = 8'hA2;
Memory[9492] = 8'h03;
Memory[9499] = 8'h00;
Memory[9498] = 8'h32;
Memory[9497] = 8'h22;
Memory[9496] = 8'hB3;
Memory[9503] = 8'h00;
Memory[9502] = 8'h02;
Memory[9501] = 8'h84;
Memory[9500] = 8'h63;
Memory[9507] = 8'h4A;
Memory[9506] = 8'h50;
Memory[9505] = 8'h50;
Memory[9504] = 8'h6F;
Memory[9511] = 8'h5F;
Memory[9510] = 8'h0C;
Memory[9509] = 8'hA2;
Memory[9508] = 8'h03;
Memory[9515] = 8'h00;
Memory[9514] = 8'h32;
Memory[9513] = 8'h22;
Memory[9512] = 8'hB3;
Memory[9519] = 8'h00;
Memory[9518] = 8'h02;
Memory[9517] = 8'h84;
Memory[9516] = 8'h63;
Memory[9523] = 8'h49;
Memory[9522] = 8'h90;
Memory[9521] = 8'h50;
Memory[9520] = 8'h6F;
Memory[9527] = 8'h5E;
Memory[9526] = 8'hCC;
Memory[9525] = 8'hA2;
Memory[9524] = 8'h03;
Memory[9531] = 8'h00;
Memory[9530] = 8'h32;
Memory[9529] = 8'h22;
Memory[9528] = 8'hB3;
Memory[9535] = 8'h00;
Memory[9534] = 8'h02;
Memory[9533] = 8'h84;
Memory[9532] = 8'h63;
Memory[9539] = 8'h48;
Memory[9538] = 8'hD0;
Memory[9537] = 8'h50;
Memory[9536] = 8'h6F;
Memory[9543] = 8'h5E;
Memory[9542] = 8'h8C;
Memory[9541] = 8'hA2;
Memory[9540] = 8'h03;
Memory[9547] = 8'h00;
Memory[9546] = 8'h32;
Memory[9545] = 8'h22;
Memory[9544] = 8'hB3;
Memory[9551] = 8'h00;
Memory[9550] = 8'h02;
Memory[9549] = 8'h84;
Memory[9548] = 8'h63;
Memory[9555] = 8'h48;
Memory[9554] = 8'h10;
Memory[9553] = 8'h50;
Memory[9552] = 8'h6F;
Memory[9559] = 8'h5E;
Memory[9558] = 8'h4C;
Memory[9557] = 8'hA2;
Memory[9556] = 8'h03;
Memory[9563] = 8'h00;
Memory[9562] = 8'h32;
Memory[9561] = 8'h22;
Memory[9560] = 8'hB3;
Memory[9567] = 8'h00;
Memory[9566] = 8'h02;
Memory[9565] = 8'h84;
Memory[9564] = 8'h63;
Memory[9571] = 8'h47;
Memory[9570] = 8'h50;
Memory[9569] = 8'h50;
Memory[9568] = 8'h6F;
Memory[9575] = 8'h5E;
Memory[9574] = 8'h0C;
Memory[9573] = 8'hA2;
Memory[9572] = 8'h03;
Memory[9579] = 8'h00;
Memory[9578] = 8'h32;
Memory[9577] = 8'h22;
Memory[9576] = 8'hB3;
Memory[9583] = 8'h00;
Memory[9582] = 8'h02;
Memory[9581] = 8'h84;
Memory[9580] = 8'h63;
Memory[9587] = 8'h46;
Memory[9586] = 8'h90;
Memory[9585] = 8'h50;
Memory[9584] = 8'h6F;
Memory[9591] = 8'h5D;
Memory[9590] = 8'hCC;
Memory[9589] = 8'hA2;
Memory[9588] = 8'h03;
Memory[9595] = 8'h00;
Memory[9594] = 8'h32;
Memory[9593] = 8'h22;
Memory[9592] = 8'hB3;
Memory[9599] = 8'h00;
Memory[9598] = 8'h02;
Memory[9597] = 8'h84;
Memory[9596] = 8'h63;
Memory[9603] = 8'h45;
Memory[9602] = 8'hD0;
Memory[9601] = 8'h50;
Memory[9600] = 8'h6F;
Memory[9607] = 8'h5D;
Memory[9606] = 8'h8C;
Memory[9605] = 8'hA2;
Memory[9604] = 8'h03;
Memory[9611] = 8'h00;
Memory[9610] = 8'h32;
Memory[9609] = 8'h22;
Memory[9608] = 8'hB3;
Memory[9615] = 8'h00;
Memory[9614] = 8'h02;
Memory[9613] = 8'h84;
Memory[9612] = 8'h63;
Memory[9619] = 8'h45;
Memory[9618] = 8'h10;
Memory[9617] = 8'h50;
Memory[9616] = 8'h6F;
Memory[9623] = 8'h5D;
Memory[9622] = 8'h4C;
Memory[9621] = 8'hA2;
Memory[9620] = 8'h03;
Memory[9627] = 8'h00;
Memory[9626] = 8'h32;
Memory[9625] = 8'h22;
Memory[9624] = 8'hB3;
Memory[9631] = 8'h00;
Memory[9630] = 8'h02;
Memory[9629] = 8'h84;
Memory[9628] = 8'h63;
Memory[9635] = 8'h44;
Memory[9634] = 8'h50;
Memory[9633] = 8'h50;
Memory[9632] = 8'h6F;
Memory[9639] = 8'h5D;
Memory[9638] = 8'h0C;
Memory[9637] = 8'hA2;
Memory[9636] = 8'h03;
Memory[9643] = 8'h00;
Memory[9642] = 8'h32;
Memory[9641] = 8'h22;
Memory[9640] = 8'hB3;
Memory[9647] = 8'h00;
Memory[9646] = 8'h02;
Memory[9645] = 8'h84;
Memory[9644] = 8'h63;
Memory[9651] = 8'h43;
Memory[9650] = 8'h90;
Memory[9649] = 8'h50;
Memory[9648] = 8'h6F;
Memory[9655] = 8'h5C;
Memory[9654] = 8'hCC;
Memory[9653] = 8'hA2;
Memory[9652] = 8'h03;
Memory[9659] = 8'h00;
Memory[9658] = 8'h32;
Memory[9657] = 8'h22;
Memory[9656] = 8'hB3;
Memory[9663] = 8'h00;
Memory[9662] = 8'h02;
Memory[9661] = 8'h84;
Memory[9660] = 8'h63;
Memory[9667] = 8'h42;
Memory[9666] = 8'hD0;
Memory[9665] = 8'h50;
Memory[9664] = 8'h6F;
Memory[9671] = 8'h5C;
Memory[9670] = 8'h8C;
Memory[9669] = 8'hA2;
Memory[9668] = 8'h03;
Memory[9675] = 8'h00;
Memory[9674] = 8'h32;
Memory[9673] = 8'h22;
Memory[9672] = 8'hB3;
Memory[9679] = 8'h00;
Memory[9678] = 8'h02;
Memory[9677] = 8'h84;
Memory[9676] = 8'h63;
Memory[9683] = 8'h42;
Memory[9682] = 8'h10;
Memory[9681] = 8'h50;
Memory[9680] = 8'h6F;
Memory[9687] = 8'h5C;
Memory[9686] = 8'h4C;
Memory[9685] = 8'hA2;
Memory[9684] = 8'h03;
Memory[9691] = 8'h00;
Memory[9690] = 8'h32;
Memory[9689] = 8'h22;
Memory[9688] = 8'hB3;
Memory[9695] = 8'h00;
Memory[9694] = 8'h02;
Memory[9693] = 8'h84;
Memory[9692] = 8'h63;
Memory[9699] = 8'h41;
Memory[9698] = 8'h50;
Memory[9697] = 8'h50;
Memory[9696] = 8'h6F;
Memory[9703] = 8'h5C;
Memory[9702] = 8'h0C;
Memory[9701] = 8'hA2;
Memory[9700] = 8'h03;
Memory[9707] = 8'h00;
Memory[9706] = 8'h32;
Memory[9705] = 8'h22;
Memory[9704] = 8'hB3;
Memory[9711] = 8'h00;
Memory[9710] = 8'h02;
Memory[9709] = 8'h84;
Memory[9708] = 8'h63;
Memory[9715] = 8'h40;
Memory[9714] = 8'h90;
Memory[9713] = 8'h50;
Memory[9712] = 8'h6F;
Memory[9719] = 8'h5B;
Memory[9718] = 8'hCC;
Memory[9717] = 8'hA2;
Memory[9716] = 8'h03;
Memory[9723] = 8'h00;
Memory[9722] = 8'h32;
Memory[9721] = 8'h22;
Memory[9720] = 8'hB3;
Memory[9727] = 8'h00;
Memory[9726] = 8'h02;
Memory[9725] = 8'h84;
Memory[9724] = 8'h63;
Memory[9731] = 8'h3F;
Memory[9730] = 8'hD0;
Memory[9729] = 8'h50;
Memory[9728] = 8'h6F;
Memory[9735] = 8'h5B;
Memory[9734] = 8'h8C;
Memory[9733] = 8'hA2;
Memory[9732] = 8'h03;
Memory[9739] = 8'h00;
Memory[9738] = 8'h32;
Memory[9737] = 8'h22;
Memory[9736] = 8'hB3;
Memory[9743] = 8'h00;
Memory[9742] = 8'h02;
Memory[9741] = 8'h84;
Memory[9740] = 8'h63;
Memory[9747] = 8'h3F;
Memory[9746] = 8'h10;
Memory[9745] = 8'h50;
Memory[9744] = 8'h6F;
Memory[9751] = 8'h5B;
Memory[9750] = 8'h4C;
Memory[9749] = 8'hA2;
Memory[9748] = 8'h03;
Memory[9755] = 8'h00;
Memory[9754] = 8'h32;
Memory[9753] = 8'h22;
Memory[9752] = 8'hB3;
Memory[9759] = 8'h00;
Memory[9758] = 8'h02;
Memory[9757] = 8'h84;
Memory[9756] = 8'h63;
Memory[9763] = 8'h3E;
Memory[9762] = 8'h50;
Memory[9761] = 8'h50;
Memory[9760] = 8'h6F;
Memory[9767] = 8'h5B;
Memory[9766] = 8'h0C;
Memory[9765] = 8'hA2;
Memory[9764] = 8'h03;
Memory[9771] = 8'h00;
Memory[9770] = 8'h32;
Memory[9769] = 8'h22;
Memory[9768] = 8'hB3;
Memory[9775] = 8'h00;
Memory[9774] = 8'h02;
Memory[9773] = 8'h84;
Memory[9772] = 8'h63;
Memory[9779] = 8'h3D;
Memory[9778] = 8'h90;
Memory[9777] = 8'h50;
Memory[9776] = 8'h6F;
Memory[9783] = 8'h5A;
Memory[9782] = 8'hCC;
Memory[9781] = 8'hA2;
Memory[9780] = 8'h03;
Memory[9787] = 8'h00;
Memory[9786] = 8'h32;
Memory[9785] = 8'h22;
Memory[9784] = 8'hB3;
Memory[9791] = 8'h00;
Memory[9790] = 8'h02;
Memory[9789] = 8'h84;
Memory[9788] = 8'h63;
Memory[9795] = 8'h3C;
Memory[9794] = 8'hD0;
Memory[9793] = 8'h50;
Memory[9792] = 8'h6F;
Memory[9799] = 8'h5A;
Memory[9798] = 8'h8C;
Memory[9797] = 8'hA2;
Memory[9796] = 8'h03;
Memory[9803] = 8'h00;
Memory[9802] = 8'h32;
Memory[9801] = 8'h22;
Memory[9800] = 8'hB3;
Memory[9807] = 8'h00;
Memory[9806] = 8'h02;
Memory[9805] = 8'h84;
Memory[9804] = 8'h63;
Memory[9811] = 8'h3C;
Memory[9810] = 8'h10;
Memory[9809] = 8'h50;
Memory[9808] = 8'h6F;
Memory[9815] = 8'h5A;
Memory[9814] = 8'h4C;
Memory[9813] = 8'hA2;
Memory[9812] = 8'h03;
Memory[9819] = 8'h00;
Memory[9818] = 8'h32;
Memory[9817] = 8'h22;
Memory[9816] = 8'hB3;
Memory[9823] = 8'h00;
Memory[9822] = 8'h02;
Memory[9821] = 8'h84;
Memory[9820] = 8'h63;
Memory[9827] = 8'h3B;
Memory[9826] = 8'h50;
Memory[9825] = 8'h50;
Memory[9824] = 8'h6F;
Memory[9831] = 8'h5A;
Memory[9830] = 8'h0C;
Memory[9829] = 8'hA2;
Memory[9828] = 8'h03;
Memory[9835] = 8'h00;
Memory[9834] = 8'h32;
Memory[9833] = 8'h22;
Memory[9832] = 8'hB3;
Memory[9839] = 8'h00;
Memory[9838] = 8'h02;
Memory[9837] = 8'h84;
Memory[9836] = 8'h63;
Memory[9843] = 8'h3A;
Memory[9842] = 8'h90;
Memory[9841] = 8'h50;
Memory[9840] = 8'h6F;
Memory[9847] = 8'h59;
Memory[9846] = 8'hCC;
Memory[9845] = 8'hA2;
Memory[9844] = 8'h03;
Memory[9851] = 8'h00;
Memory[9850] = 8'h32;
Memory[9849] = 8'h22;
Memory[9848] = 8'hB3;
Memory[9855] = 8'h00;
Memory[9854] = 8'h02;
Memory[9853] = 8'h84;
Memory[9852] = 8'h63;
Memory[9859] = 8'h39;
Memory[9858] = 8'hD0;
Memory[9857] = 8'h50;
Memory[9856] = 8'h6F;
Memory[9863] = 8'h59;
Memory[9862] = 8'h8C;
Memory[9861] = 8'hA2;
Memory[9860] = 8'h03;
Memory[9867] = 8'h00;
Memory[9866] = 8'h32;
Memory[9865] = 8'h22;
Memory[9864] = 8'hB3;
Memory[9871] = 8'h00;
Memory[9870] = 8'h02;
Memory[9869] = 8'h84;
Memory[9868] = 8'h63;
Memory[9875] = 8'h39;
Memory[9874] = 8'h10;
Memory[9873] = 8'h50;
Memory[9872] = 8'h6F;
Memory[9879] = 8'h59;
Memory[9878] = 8'h4C;
Memory[9877] = 8'hA2;
Memory[9876] = 8'h03;
Memory[9883] = 8'h00;
Memory[9882] = 8'h32;
Memory[9881] = 8'h22;
Memory[9880] = 8'hB3;
Memory[9887] = 8'h00;
Memory[9886] = 8'h02;
Memory[9885] = 8'h84;
Memory[9884] = 8'h63;
Memory[9891] = 8'h38;
Memory[9890] = 8'h50;
Memory[9889] = 8'h50;
Memory[9888] = 8'h6F;
Memory[9895] = 8'h59;
Memory[9894] = 8'h0C;
Memory[9893] = 8'hA2;
Memory[9892] = 8'h03;
Memory[9899] = 8'h00;
Memory[9898] = 8'h32;
Memory[9897] = 8'h22;
Memory[9896] = 8'hB3;
Memory[9903] = 8'h00;
Memory[9902] = 8'h02;
Memory[9901] = 8'h84;
Memory[9900] = 8'h63;
Memory[9907] = 8'h37;
Memory[9906] = 8'h90;
Memory[9905] = 8'h50;
Memory[9904] = 8'h6F;
Memory[9911] = 8'h58;
Memory[9910] = 8'hCC;
Memory[9909] = 8'hA2;
Memory[9908] = 8'h03;
Memory[9915] = 8'h00;
Memory[9914] = 8'h32;
Memory[9913] = 8'h22;
Memory[9912] = 8'hB3;
Memory[9919] = 8'h00;
Memory[9918] = 8'h02;
Memory[9917] = 8'h84;
Memory[9916] = 8'h63;
Memory[9923] = 8'h36;
Memory[9922] = 8'hD0;
Memory[9921] = 8'h50;
Memory[9920] = 8'h6F;
Memory[9927] = 8'h58;
Memory[9926] = 8'h8C;
Memory[9925] = 8'hA2;
Memory[9924] = 8'h03;
Memory[9931] = 8'h00;
Memory[9930] = 8'h32;
Memory[9929] = 8'h22;
Memory[9928] = 8'hB3;
Memory[9935] = 8'h00;
Memory[9934] = 8'h02;
Memory[9933] = 8'h84;
Memory[9932] = 8'h63;
Memory[9939] = 8'h36;
Memory[9938] = 8'h10;
Memory[9937] = 8'h50;
Memory[9936] = 8'h6F;
Memory[9943] = 8'h58;
Memory[9942] = 8'h4C;
Memory[9941] = 8'hA2;
Memory[9940] = 8'h03;
Memory[9947] = 8'h00;
Memory[9946] = 8'h32;
Memory[9945] = 8'h22;
Memory[9944] = 8'hB3;
Memory[9951] = 8'h00;
Memory[9950] = 8'h02;
Memory[9949] = 8'h84;
Memory[9948] = 8'h63;
Memory[9955] = 8'h35;
Memory[9954] = 8'h50;
Memory[9953] = 8'h50;
Memory[9952] = 8'h6F;
Memory[9959] = 8'h58;
Memory[9958] = 8'h0C;
Memory[9957] = 8'hA2;
Memory[9956] = 8'h03;
Memory[9963] = 8'h00;
Memory[9962] = 8'h32;
Memory[9961] = 8'h22;
Memory[9960] = 8'hB3;
Memory[9967] = 8'h00;
Memory[9966] = 8'h02;
Memory[9965] = 8'h84;
Memory[9964] = 8'h63;
Memory[9971] = 8'h34;
Memory[9970] = 8'h90;
Memory[9969] = 8'h50;
Memory[9968] = 8'h6F;
Memory[9975] = 8'h57;
Memory[9974] = 8'hCC;
Memory[9973] = 8'hA2;
Memory[9972] = 8'h03;
Memory[9979] = 8'h00;
Memory[9978] = 8'h32;
Memory[9977] = 8'h22;
Memory[9976] = 8'hB3;
Memory[9983] = 8'h00;
Memory[9982] = 8'h02;
Memory[9981] = 8'h84;
Memory[9980] = 8'h63;
Memory[9987] = 8'h33;
Memory[9986] = 8'hD0;
Memory[9985] = 8'h50;
Memory[9984] = 8'h6F;
Memory[9991] = 8'h57;
Memory[9990] = 8'h8C;
Memory[9989] = 8'hA2;
Memory[9988] = 8'h03;
Memory[9995] = 8'h00;
Memory[9994] = 8'h32;
Memory[9993] = 8'h22;
Memory[9992] = 8'hB3;
Memory[9999] = 8'h00;
Memory[9998] = 8'h02;
Memory[9997] = 8'h84;
Memory[9996] = 8'h63;
Memory[10003] = 8'h33;
Memory[10002] = 8'h10;
Memory[10001] = 8'h50;
Memory[10000] = 8'h6F;
Memory[10007] = 8'h57;
Memory[10006] = 8'h4C;
Memory[10005] = 8'hA2;
Memory[10004] = 8'h03;
Memory[10011] = 8'h00;
Memory[10010] = 8'h32;
Memory[10009] = 8'h22;
Memory[10008] = 8'hB3;
Memory[10015] = 8'h00;
Memory[10014] = 8'h02;
Memory[10013] = 8'h84;
Memory[10012] = 8'h63;
Memory[10019] = 8'h32;
Memory[10018] = 8'h50;
Memory[10017] = 8'h50;
Memory[10016] = 8'h6F;
Memory[10023] = 8'h57;
Memory[10022] = 8'h0C;
Memory[10021] = 8'hA2;
Memory[10020] = 8'h03;
Memory[10027] = 8'h00;
Memory[10026] = 8'h32;
Memory[10025] = 8'h22;
Memory[10024] = 8'hB3;
Memory[10031] = 8'h00;
Memory[10030] = 8'h02;
Memory[10029] = 8'h84;
Memory[10028] = 8'h63;
Memory[10035] = 8'h31;
Memory[10034] = 8'h90;
Memory[10033] = 8'h50;
Memory[10032] = 8'h6F;
Memory[10039] = 8'h56;
Memory[10038] = 8'hCC;
Memory[10037] = 8'hA2;
Memory[10036] = 8'h03;
Memory[10043] = 8'h00;
Memory[10042] = 8'h32;
Memory[10041] = 8'h22;
Memory[10040] = 8'hB3;
Memory[10047] = 8'h00;
Memory[10046] = 8'h02;
Memory[10045] = 8'h84;
Memory[10044] = 8'h63;
Memory[10051] = 8'h30;
Memory[10050] = 8'hD0;
Memory[10049] = 8'h50;
Memory[10048] = 8'h6F;
Memory[10055] = 8'h56;
Memory[10054] = 8'h8C;
Memory[10053] = 8'hA2;
Memory[10052] = 8'h03;
Memory[10059] = 8'h00;
Memory[10058] = 8'h32;
Memory[10057] = 8'h22;
Memory[10056] = 8'hB3;
Memory[10063] = 8'h00;
Memory[10062] = 8'h02;
Memory[10061] = 8'h84;
Memory[10060] = 8'h63;
Memory[10067] = 8'h30;
Memory[10066] = 8'h10;
Memory[10065] = 8'h50;
Memory[10064] = 8'h6F;
Memory[10071] = 8'h56;
Memory[10070] = 8'h4C;
Memory[10069] = 8'hA2;
Memory[10068] = 8'h03;
Memory[10075] = 8'h00;
Memory[10074] = 8'h32;
Memory[10073] = 8'h22;
Memory[10072] = 8'hB3;
Memory[10079] = 8'h00;
Memory[10078] = 8'h02;
Memory[10077] = 8'h84;
Memory[10076] = 8'h63;
Memory[10083] = 8'h2F;
Memory[10082] = 8'h50;
Memory[10081] = 8'h50;
Memory[10080] = 8'h6F;
Memory[10087] = 8'h56;
Memory[10086] = 8'h0C;
Memory[10085] = 8'hA2;
Memory[10084] = 8'h03;
Memory[10091] = 8'h00;
Memory[10090] = 8'h32;
Memory[10089] = 8'h22;
Memory[10088] = 8'hB3;
Memory[10095] = 8'h00;
Memory[10094] = 8'h02;
Memory[10093] = 8'h84;
Memory[10092] = 8'h63;
Memory[10099] = 8'h2E;
Memory[10098] = 8'h90;
Memory[10097] = 8'h50;
Memory[10096] = 8'h6F;
Memory[10103] = 8'h55;
Memory[10102] = 8'hCC;
Memory[10101] = 8'hA2;
Memory[10100] = 8'h03;
Memory[10107] = 8'h00;
Memory[10106] = 8'h32;
Memory[10105] = 8'h22;
Memory[10104] = 8'hB3;
Memory[10111] = 8'h00;
Memory[10110] = 8'h02;
Memory[10109] = 8'h84;
Memory[10108] = 8'h63;
Memory[10115] = 8'h2D;
Memory[10114] = 8'hD0;
Memory[10113] = 8'h50;
Memory[10112] = 8'h6F;
Memory[10119] = 8'h55;
Memory[10118] = 8'h8C;
Memory[10117] = 8'hA2;
Memory[10116] = 8'h03;
Memory[10123] = 8'h00;
Memory[10122] = 8'h32;
Memory[10121] = 8'h22;
Memory[10120] = 8'hB3;
Memory[10127] = 8'h00;
Memory[10126] = 8'h02;
Memory[10125] = 8'h84;
Memory[10124] = 8'h63;
Memory[10131] = 8'h2D;
Memory[10130] = 8'h10;
Memory[10129] = 8'h50;
Memory[10128] = 8'h6F;
Memory[10135] = 8'h55;
Memory[10134] = 8'h4C;
Memory[10133] = 8'hA2;
Memory[10132] = 8'h03;
Memory[10139] = 8'h00;
Memory[10138] = 8'h32;
Memory[10137] = 8'h22;
Memory[10136] = 8'hB3;
Memory[10143] = 8'h00;
Memory[10142] = 8'h02;
Memory[10141] = 8'h84;
Memory[10140] = 8'h63;
Memory[10147] = 8'h2C;
Memory[10146] = 8'h50;
Memory[10145] = 8'h50;
Memory[10144] = 8'h6F;
Memory[10151] = 8'h55;
Memory[10150] = 8'h0C;
Memory[10149] = 8'hA2;
Memory[10148] = 8'h03;
Memory[10155] = 8'h00;
Memory[10154] = 8'h32;
Memory[10153] = 8'h22;
Memory[10152] = 8'hB3;
Memory[10159] = 8'h00;
Memory[10158] = 8'h02;
Memory[10157] = 8'h84;
Memory[10156] = 8'h63;
Memory[10163] = 8'h2B;
Memory[10162] = 8'h90;
Memory[10161] = 8'h50;
Memory[10160] = 8'h6F;
Memory[10167] = 8'h54;
Memory[10166] = 8'hCC;
Memory[10165] = 8'hA2;
Memory[10164] = 8'h03;
Memory[10171] = 8'h00;
Memory[10170] = 8'h32;
Memory[10169] = 8'h22;
Memory[10168] = 8'hB3;
Memory[10175] = 8'h00;
Memory[10174] = 8'h02;
Memory[10173] = 8'h84;
Memory[10172] = 8'h63;
Memory[10179] = 8'h2A;
Memory[10178] = 8'hD0;
Memory[10177] = 8'h50;
Memory[10176] = 8'h6F;
Memory[10183] = 8'h54;
Memory[10182] = 8'h8C;
Memory[10181] = 8'hA2;
Memory[10180] = 8'h03;
Memory[10187] = 8'h00;
Memory[10186] = 8'h32;
Memory[10185] = 8'h22;
Memory[10184] = 8'hB3;
Memory[10191] = 8'h00;
Memory[10190] = 8'h02;
Memory[10189] = 8'h84;
Memory[10188] = 8'h63;
Memory[10195] = 8'h2A;
Memory[10194] = 8'h10;
Memory[10193] = 8'h50;
Memory[10192] = 8'h6F;
Memory[10199] = 8'h54;
Memory[10198] = 8'h4C;
Memory[10197] = 8'hA2;
Memory[10196] = 8'h03;
Memory[10203] = 8'h00;
Memory[10202] = 8'h32;
Memory[10201] = 8'h22;
Memory[10200] = 8'hB3;
Memory[10207] = 8'h00;
Memory[10206] = 8'h02;
Memory[10205] = 8'h84;
Memory[10204] = 8'h63;
Memory[10211] = 8'h29;
Memory[10210] = 8'h50;
Memory[10209] = 8'h50;
Memory[10208] = 8'h6F;
Memory[10215] = 8'h54;
Memory[10214] = 8'h0C;
Memory[10213] = 8'hA2;
Memory[10212] = 8'h03;
Memory[10219] = 8'h00;
Memory[10218] = 8'h32;
Memory[10217] = 8'h22;
Memory[10216] = 8'hB3;
Memory[10223] = 8'h00;
Memory[10222] = 8'h02;
Memory[10221] = 8'h84;
Memory[10220] = 8'h63;
Memory[10227] = 8'h28;
Memory[10226] = 8'h90;
Memory[10225] = 8'h50;
Memory[10224] = 8'h6F;
Memory[10231] = 8'h53;
Memory[10230] = 8'hCC;
Memory[10229] = 8'hA2;
Memory[10228] = 8'h03;
Memory[10235] = 8'h00;
Memory[10234] = 8'h32;
Memory[10233] = 8'h22;
Memory[10232] = 8'hB3;
Memory[10239] = 8'h00;
Memory[10238] = 8'h02;
Memory[10237] = 8'h84;
Memory[10236] = 8'h63;
Memory[10243] = 8'h27;
Memory[10242] = 8'hD0;
Memory[10241] = 8'h50;
Memory[10240] = 8'h6F;
Memory[10247] = 8'h53;
Memory[10246] = 8'h8C;
Memory[10245] = 8'hA2;
Memory[10244] = 8'h03;
Memory[10251] = 8'h00;
Memory[10250] = 8'h32;
Memory[10249] = 8'h22;
Memory[10248] = 8'hB3;
Memory[10255] = 8'h00;
Memory[10254] = 8'h02;
Memory[10253] = 8'h84;
Memory[10252] = 8'h63;
Memory[10259] = 8'h27;
Memory[10258] = 8'h10;
Memory[10257] = 8'h50;
Memory[10256] = 8'h6F;
Memory[10263] = 8'h53;
Memory[10262] = 8'h4C;
Memory[10261] = 8'hA2;
Memory[10260] = 8'h03;
Memory[10267] = 8'h00;
Memory[10266] = 8'h32;
Memory[10265] = 8'h22;
Memory[10264] = 8'hB3;
Memory[10271] = 8'h00;
Memory[10270] = 8'h02;
Memory[10269] = 8'h84;
Memory[10268] = 8'h63;
Memory[10275] = 8'h26;
Memory[10274] = 8'h50;
Memory[10273] = 8'h50;
Memory[10272] = 8'h6F;
Memory[10279] = 8'h53;
Memory[10278] = 8'h0C;
Memory[10277] = 8'hA2;
Memory[10276] = 8'h03;
Memory[10283] = 8'h00;
Memory[10282] = 8'h32;
Memory[10281] = 8'h22;
Memory[10280] = 8'hB3;
Memory[10287] = 8'h00;
Memory[10286] = 8'h02;
Memory[10285] = 8'h84;
Memory[10284] = 8'h63;
Memory[10291] = 8'h25;
Memory[10290] = 8'h90;
Memory[10289] = 8'h50;
Memory[10288] = 8'h6F;
Memory[10295] = 8'h52;
Memory[10294] = 8'hCC;
Memory[10293] = 8'hA2;
Memory[10292] = 8'h03;
Memory[10299] = 8'h00;
Memory[10298] = 8'h32;
Memory[10297] = 8'h22;
Memory[10296] = 8'hB3;
Memory[10303] = 8'h00;
Memory[10302] = 8'h02;
Memory[10301] = 8'h84;
Memory[10300] = 8'h63;
Memory[10307] = 8'h24;
Memory[10306] = 8'hD0;
Memory[10305] = 8'h50;
Memory[10304] = 8'h6F;
Memory[10311] = 8'h52;
Memory[10310] = 8'h8C;
Memory[10309] = 8'hA2;
Memory[10308] = 8'h03;
Memory[10315] = 8'h00;
Memory[10314] = 8'h32;
Memory[10313] = 8'h22;
Memory[10312] = 8'hB3;
Memory[10319] = 8'h00;
Memory[10318] = 8'h02;
Memory[10317] = 8'h84;
Memory[10316] = 8'h63;
Memory[10323] = 8'h24;
Memory[10322] = 8'h10;
Memory[10321] = 8'h50;
Memory[10320] = 8'h6F;
Memory[10327] = 8'h52;
Memory[10326] = 8'h4C;
Memory[10325] = 8'hA2;
Memory[10324] = 8'h03;
Memory[10331] = 8'h00;
Memory[10330] = 8'h32;
Memory[10329] = 8'h22;
Memory[10328] = 8'hB3;
Memory[10335] = 8'h00;
Memory[10334] = 8'h02;
Memory[10333] = 8'h84;
Memory[10332] = 8'h63;
Memory[10339] = 8'h23;
Memory[10338] = 8'h50;
Memory[10337] = 8'h50;
Memory[10336] = 8'h6F;
Memory[10343] = 8'h52;
Memory[10342] = 8'h0C;
Memory[10341] = 8'hA2;
Memory[10340] = 8'h03;
Memory[10347] = 8'h00;
Memory[10346] = 8'h32;
Memory[10345] = 8'h22;
Memory[10344] = 8'hB3;
Memory[10351] = 8'h00;
Memory[10350] = 8'h02;
Memory[10349] = 8'h84;
Memory[10348] = 8'h63;
Memory[10355] = 8'h22;
Memory[10354] = 8'h90;
Memory[10353] = 8'h50;
Memory[10352] = 8'h6F;
Memory[10359] = 8'h51;
Memory[10358] = 8'hCC;
Memory[10357] = 8'hA2;
Memory[10356] = 8'h03;
Memory[10363] = 8'h00;
Memory[10362] = 8'h32;
Memory[10361] = 8'h22;
Memory[10360] = 8'hB3;
Memory[10367] = 8'h00;
Memory[10366] = 8'h02;
Memory[10365] = 8'h84;
Memory[10364] = 8'h63;
Memory[10371] = 8'h21;
Memory[10370] = 8'hD0;
Memory[10369] = 8'h50;
Memory[10368] = 8'h6F;
Memory[10375] = 8'h51;
Memory[10374] = 8'h8C;
Memory[10373] = 8'hA2;
Memory[10372] = 8'h03;
Memory[10379] = 8'h00;
Memory[10378] = 8'h32;
Memory[10377] = 8'h22;
Memory[10376] = 8'hB3;
Memory[10383] = 8'h00;
Memory[10382] = 8'h02;
Memory[10381] = 8'h84;
Memory[10380] = 8'h63;
Memory[10387] = 8'h21;
Memory[10386] = 8'h10;
Memory[10385] = 8'h50;
Memory[10384] = 8'h6F;
Memory[10391] = 8'h51;
Memory[10390] = 8'h4C;
Memory[10389] = 8'hA2;
Memory[10388] = 8'h03;
Memory[10395] = 8'h00;
Memory[10394] = 8'h32;
Memory[10393] = 8'h22;
Memory[10392] = 8'hB3;
Memory[10399] = 8'h00;
Memory[10398] = 8'h02;
Memory[10397] = 8'h84;
Memory[10396] = 8'h63;
Memory[10403] = 8'h20;
Memory[10402] = 8'h50;
Memory[10401] = 8'h50;
Memory[10400] = 8'h6F;
Memory[10407] = 8'h51;
Memory[10406] = 8'h0C;
Memory[10405] = 8'hA2;
Memory[10404] = 8'h03;
Memory[10411] = 8'h00;
Memory[10410] = 8'h32;
Memory[10409] = 8'h22;
Memory[10408] = 8'hB3;
Memory[10415] = 8'h00;
Memory[10414] = 8'h02;
Memory[10413] = 8'h84;
Memory[10412] = 8'h63;
Memory[10419] = 8'h1F;
Memory[10418] = 8'h90;
Memory[10417] = 8'h50;
Memory[10416] = 8'h6F;
Memory[10423] = 8'h50;
Memory[10422] = 8'hCC;
Memory[10421] = 8'hA2;
Memory[10420] = 8'h03;
Memory[10427] = 8'h00;
Memory[10426] = 8'h32;
Memory[10425] = 8'h22;
Memory[10424] = 8'hB3;
Memory[10431] = 8'h00;
Memory[10430] = 8'h02;
Memory[10429] = 8'h84;
Memory[10428] = 8'h63;
Memory[10435] = 8'h1E;
Memory[10434] = 8'hD0;
Memory[10433] = 8'h50;
Memory[10432] = 8'h6F;
Memory[10439] = 8'h50;
Memory[10438] = 8'h8C;
Memory[10437] = 8'hA2;
Memory[10436] = 8'h03;
Memory[10443] = 8'h00;
Memory[10442] = 8'h32;
Memory[10441] = 8'h22;
Memory[10440] = 8'hB3;
Memory[10447] = 8'h00;
Memory[10446] = 8'h02;
Memory[10445] = 8'h84;
Memory[10444] = 8'h63;
Memory[10451] = 8'h1E;
Memory[10450] = 8'h10;
Memory[10449] = 8'h50;
Memory[10448] = 8'h6F;
Memory[10455] = 8'h50;
Memory[10454] = 8'h4C;
Memory[10453] = 8'hA2;
Memory[10452] = 8'h03;
Memory[10459] = 8'h00;
Memory[10458] = 8'h32;
Memory[10457] = 8'h22;
Memory[10456] = 8'hB3;
Memory[10463] = 8'h00;
Memory[10462] = 8'h02;
Memory[10461] = 8'h84;
Memory[10460] = 8'h63;
Memory[10467] = 8'h1D;
Memory[10466] = 8'h50;
Memory[10465] = 8'h50;
Memory[10464] = 8'h6F;
Memory[10471] = 8'h50;
Memory[10470] = 8'h0C;
Memory[10469] = 8'hA2;
Memory[10468] = 8'h03;
Memory[10475] = 8'h00;
Memory[10474] = 8'h32;
Memory[10473] = 8'h22;
Memory[10472] = 8'hB3;
Memory[10479] = 8'h00;
Memory[10478] = 8'h02;
Memory[10477] = 8'h84;
Memory[10476] = 8'h63;
Memory[10483] = 8'h1C;
Memory[10482] = 8'h90;
Memory[10481] = 8'h50;
Memory[10480] = 8'h6F;
Memory[10487] = 8'h4F;
Memory[10486] = 8'hCC;
Memory[10485] = 8'hA2;
Memory[10484] = 8'h03;
Memory[10491] = 8'h00;
Memory[10490] = 8'h32;
Memory[10489] = 8'h22;
Memory[10488] = 8'hB3;
Memory[10495] = 8'h00;
Memory[10494] = 8'h02;
Memory[10493] = 8'h84;
Memory[10492] = 8'h63;
Memory[10499] = 8'h1B;
Memory[10498] = 8'hD0;
Memory[10497] = 8'h50;
Memory[10496] = 8'h6F;
Memory[10503] = 8'h4F;
Memory[10502] = 8'h8C;
Memory[10501] = 8'hA2;
Memory[10500] = 8'h03;
Memory[10507] = 8'h00;
Memory[10506] = 8'h32;
Memory[10505] = 8'h22;
Memory[10504] = 8'hB3;
Memory[10511] = 8'h00;
Memory[10510] = 8'h02;
Memory[10509] = 8'h84;
Memory[10508] = 8'h63;
Memory[10515] = 8'h1B;
Memory[10514] = 8'h10;
Memory[10513] = 8'h50;
Memory[10512] = 8'h6F;
Memory[10519] = 8'h4F;
Memory[10518] = 8'h4C;
Memory[10517] = 8'hA2;
Memory[10516] = 8'h03;
Memory[10523] = 8'h00;
Memory[10522] = 8'h32;
Memory[10521] = 8'h22;
Memory[10520] = 8'hB3;
Memory[10527] = 8'h00;
Memory[10526] = 8'h02;
Memory[10525] = 8'h84;
Memory[10524] = 8'h63;
Memory[10531] = 8'h1A;
Memory[10530] = 8'h50;
Memory[10529] = 8'h50;
Memory[10528] = 8'h6F;
Memory[10535] = 8'h4F;
Memory[10534] = 8'h0C;
Memory[10533] = 8'hA2;
Memory[10532] = 8'h03;
Memory[10539] = 8'h00;
Memory[10538] = 8'h32;
Memory[10537] = 8'h22;
Memory[10536] = 8'hB3;
Memory[10543] = 8'h00;
Memory[10542] = 8'h02;
Memory[10541] = 8'h84;
Memory[10540] = 8'h63;
Memory[10547] = 8'h19;
Memory[10546] = 8'h90;
Memory[10545] = 8'h50;
Memory[10544] = 8'h6F;
Memory[10551] = 8'h4E;
Memory[10550] = 8'hCC;
Memory[10549] = 8'hA2;
Memory[10548] = 8'h03;
Memory[10555] = 8'h00;
Memory[10554] = 8'h32;
Memory[10553] = 8'h22;
Memory[10552] = 8'hB3;
Memory[10559] = 8'h00;
Memory[10558] = 8'h02;
Memory[10557] = 8'h84;
Memory[10556] = 8'h63;
Memory[10563] = 8'h18;
Memory[10562] = 8'hD0;
Memory[10561] = 8'h50;
Memory[10560] = 8'h6F;
Memory[10567] = 8'h4E;
Memory[10566] = 8'h8C;
Memory[10565] = 8'hA2;
Memory[10564] = 8'h03;
Memory[10571] = 8'h00;
Memory[10570] = 8'h32;
Memory[10569] = 8'h22;
Memory[10568] = 8'hB3;
Memory[10575] = 8'h00;
Memory[10574] = 8'h02;
Memory[10573] = 8'h84;
Memory[10572] = 8'h63;
Memory[10579] = 8'h18;
Memory[10578] = 8'h10;
Memory[10577] = 8'h50;
Memory[10576] = 8'h6F;
Memory[10583] = 8'h4E;
Memory[10582] = 8'h4C;
Memory[10581] = 8'hA2;
Memory[10580] = 8'h03;
Memory[10587] = 8'h00;
Memory[10586] = 8'h32;
Memory[10585] = 8'h22;
Memory[10584] = 8'hB3;
Memory[10591] = 8'h00;
Memory[10590] = 8'h02;
Memory[10589] = 8'h84;
Memory[10588] = 8'h63;
Memory[10595] = 8'h17;
Memory[10594] = 8'h50;
Memory[10593] = 8'h50;
Memory[10592] = 8'h6F;
Memory[10599] = 8'h4E;
Memory[10598] = 8'h0C;
Memory[10597] = 8'hA2;
Memory[10596] = 8'h03;
Memory[10603] = 8'h00;
Memory[10602] = 8'h32;
Memory[10601] = 8'h22;
Memory[10600] = 8'hB3;
Memory[10607] = 8'h00;
Memory[10606] = 8'h02;
Memory[10605] = 8'h84;
Memory[10604] = 8'h63;
Memory[10611] = 8'h16;
Memory[10610] = 8'h90;
Memory[10609] = 8'h50;
Memory[10608] = 8'h6F;
Memory[10615] = 8'h4D;
Memory[10614] = 8'hCC;
Memory[10613] = 8'hA2;
Memory[10612] = 8'h03;
Memory[10619] = 8'h00;
Memory[10618] = 8'h32;
Memory[10617] = 8'h22;
Memory[10616] = 8'hB3;
Memory[10623] = 8'h00;
Memory[10622] = 8'h02;
Memory[10621] = 8'h84;
Memory[10620] = 8'h63;
Memory[10627] = 8'h15;
Memory[10626] = 8'hD0;
Memory[10625] = 8'h50;
Memory[10624] = 8'h6F;
Memory[10631] = 8'h4D;
Memory[10630] = 8'h8C;
Memory[10629] = 8'hA2;
Memory[10628] = 8'h03;
Memory[10635] = 8'h00;
Memory[10634] = 8'h32;
Memory[10633] = 8'h22;
Memory[10632] = 8'hB3;
Memory[10639] = 8'h00;
Memory[10638] = 8'h02;
Memory[10637] = 8'h84;
Memory[10636] = 8'h63;
Memory[10643] = 8'h15;
Memory[10642] = 8'h10;
Memory[10641] = 8'h50;
Memory[10640] = 8'h6F;
Memory[10647] = 8'h4D;
Memory[10646] = 8'h4C;
Memory[10645] = 8'hA2;
Memory[10644] = 8'h03;
Memory[10651] = 8'h00;
Memory[10650] = 8'h32;
Memory[10649] = 8'h22;
Memory[10648] = 8'hB3;
Memory[10655] = 8'h00;
Memory[10654] = 8'h02;
Memory[10653] = 8'h84;
Memory[10652] = 8'h63;
Memory[10659] = 8'h14;
Memory[10658] = 8'h50;
Memory[10657] = 8'h50;
Memory[10656] = 8'h6F;
Memory[10663] = 8'h4D;
Memory[10662] = 8'h0C;
Memory[10661] = 8'hA2;
Memory[10660] = 8'h03;
Memory[10667] = 8'h00;
Memory[10666] = 8'h32;
Memory[10665] = 8'h22;
Memory[10664] = 8'hB3;
Memory[10671] = 8'h00;
Memory[10670] = 8'h02;
Memory[10669] = 8'h84;
Memory[10668] = 8'h63;
Memory[10675] = 8'h13;
Memory[10674] = 8'h90;
Memory[10673] = 8'h50;
Memory[10672] = 8'h6F;
Memory[10679] = 8'h4C;
Memory[10678] = 8'hCC;
Memory[10677] = 8'hA2;
Memory[10676] = 8'h03;
Memory[10683] = 8'h00;
Memory[10682] = 8'h32;
Memory[10681] = 8'h22;
Memory[10680] = 8'hB3;
Memory[10687] = 8'h00;
Memory[10686] = 8'h02;
Memory[10685] = 8'h84;
Memory[10684] = 8'h63;
Memory[10691] = 8'h12;
Memory[10690] = 8'hD0;
Memory[10689] = 8'h50;
Memory[10688] = 8'h6F;
Memory[10695] = 8'h4C;
Memory[10694] = 8'h8C;
Memory[10693] = 8'hA2;
Memory[10692] = 8'h03;
Memory[10699] = 8'h00;
Memory[10698] = 8'h32;
Memory[10697] = 8'h22;
Memory[10696] = 8'hB3;
Memory[10703] = 8'h00;
Memory[10702] = 8'h02;
Memory[10701] = 8'h84;
Memory[10700] = 8'h63;
Memory[10707] = 8'h12;
Memory[10706] = 8'h10;
Memory[10705] = 8'h50;
Memory[10704] = 8'h6F;
Memory[10711] = 8'h4C;
Memory[10710] = 8'h4C;
Memory[10709] = 8'hA2;
Memory[10708] = 8'h03;
Memory[10715] = 8'h00;
Memory[10714] = 8'h32;
Memory[10713] = 8'h22;
Memory[10712] = 8'hB3;
Memory[10719] = 8'h00;
Memory[10718] = 8'h02;
Memory[10717] = 8'h84;
Memory[10716] = 8'h63;
Memory[10723] = 8'h11;
Memory[10722] = 8'h50;
Memory[10721] = 8'h50;
Memory[10720] = 8'h6F;
Memory[10727] = 8'h4C;
Memory[10726] = 8'h0C;
Memory[10725] = 8'hA2;
Memory[10724] = 8'h03;
Memory[10731] = 8'h00;
Memory[10730] = 8'h32;
Memory[10729] = 8'h22;
Memory[10728] = 8'hB3;
Memory[10735] = 8'h00;
Memory[10734] = 8'h02;
Memory[10733] = 8'h84;
Memory[10732] = 8'h63;
Memory[10739] = 8'h10;
Memory[10738] = 8'h90;
Memory[10737] = 8'h50;
Memory[10736] = 8'h6F;
Memory[10743] = 8'h4B;
Memory[10742] = 8'hCC;
Memory[10741] = 8'hA2;
Memory[10740] = 8'h03;
Memory[10747] = 8'h00;
Memory[10746] = 8'h32;
Memory[10745] = 8'h22;
Memory[10744] = 8'hB3;
Memory[10751] = 8'h00;
Memory[10750] = 8'h02;
Memory[10749] = 8'h84;
Memory[10748] = 8'h63;
Memory[10755] = 8'h0F;
Memory[10754] = 8'hD0;
Memory[10753] = 8'h50;
Memory[10752] = 8'h6F;
Memory[10759] = 8'h4B;
Memory[10758] = 8'h8C;
Memory[10757] = 8'hA2;
Memory[10756] = 8'h03;
Memory[10763] = 8'h00;
Memory[10762] = 8'h32;
Memory[10761] = 8'h22;
Memory[10760] = 8'hB3;
Memory[10767] = 8'h00;
Memory[10766] = 8'h02;
Memory[10765] = 8'h84;
Memory[10764] = 8'h63;
Memory[10771] = 8'h0F;
Memory[10770] = 8'h10;
Memory[10769] = 8'h50;
Memory[10768] = 8'h6F;
Memory[10775] = 8'h4B;
Memory[10774] = 8'h4C;
Memory[10773] = 8'hA2;
Memory[10772] = 8'h03;
Memory[10779] = 8'h00;
Memory[10778] = 8'h32;
Memory[10777] = 8'h22;
Memory[10776] = 8'hB3;
Memory[10783] = 8'h00;
Memory[10782] = 8'h02;
Memory[10781] = 8'h84;
Memory[10780] = 8'h63;
Memory[10787] = 8'h0E;
Memory[10786] = 8'h50;
Memory[10785] = 8'h50;
Memory[10784] = 8'h6F;
Memory[10791] = 8'h4B;
Memory[10790] = 8'h0C;
Memory[10789] = 8'hA2;
Memory[10788] = 8'h03;
Memory[10795] = 8'h00;
Memory[10794] = 8'h32;
Memory[10793] = 8'h22;
Memory[10792] = 8'hB3;
Memory[10799] = 8'h00;
Memory[10798] = 8'h02;
Memory[10797] = 8'h84;
Memory[10796] = 8'h63;
Memory[10803] = 8'h0D;
Memory[10802] = 8'h90;
Memory[10801] = 8'h50;
Memory[10800] = 8'h6F;
Memory[10807] = 8'h4A;
Memory[10806] = 8'hCC;
Memory[10805] = 8'hA2;
Memory[10804] = 8'h03;
Memory[10811] = 8'h00;
Memory[10810] = 8'h32;
Memory[10809] = 8'h22;
Memory[10808] = 8'hB3;
Memory[10815] = 8'h00;
Memory[10814] = 8'h02;
Memory[10813] = 8'h84;
Memory[10812] = 8'h63;
Memory[10819] = 8'h0C;
Memory[10818] = 8'hD0;
Memory[10817] = 8'h50;
Memory[10816] = 8'h6F;
Memory[10823] = 8'h4A;
Memory[10822] = 8'h8C;
Memory[10821] = 8'hA2;
Memory[10820] = 8'h03;
Memory[10827] = 8'h00;
Memory[10826] = 8'h32;
Memory[10825] = 8'h22;
Memory[10824] = 8'hB3;
Memory[10831] = 8'h00;
Memory[10830] = 8'h02;
Memory[10829] = 8'h84;
Memory[10828] = 8'h63;
Memory[10835] = 8'h0C;
Memory[10834] = 8'h10;
Memory[10833] = 8'h50;
Memory[10832] = 8'h6F;
Memory[10839] = 8'h4A;
Memory[10838] = 8'h4C;
Memory[10837] = 8'hA2;
Memory[10836] = 8'h03;
Memory[10843] = 8'h00;
Memory[10842] = 8'h32;
Memory[10841] = 8'h22;
Memory[10840] = 8'hB3;
Memory[10847] = 8'h00;
Memory[10846] = 8'h02;
Memory[10845] = 8'h84;
Memory[10844] = 8'h63;
Memory[10851] = 8'h0B;
Memory[10850] = 8'h50;
Memory[10849] = 8'h50;
Memory[10848] = 8'h6F;
Memory[10855] = 8'h4A;
Memory[10854] = 8'h0C;
Memory[10853] = 8'hA2;
Memory[10852] = 8'h03;
Memory[10859] = 8'h00;
Memory[10858] = 8'h32;
Memory[10857] = 8'h22;
Memory[10856] = 8'hB3;
Memory[10863] = 8'h00;
Memory[10862] = 8'h02;
Memory[10861] = 8'h84;
Memory[10860] = 8'h63;
Memory[10867] = 8'h0A;
Memory[10866] = 8'h90;
Memory[10865] = 8'h50;
Memory[10864] = 8'h6F;
Memory[10871] = 8'h49;
Memory[10870] = 8'hCC;
Memory[10869] = 8'hA2;
Memory[10868] = 8'h03;
Memory[10875] = 8'h00;
Memory[10874] = 8'h32;
Memory[10873] = 8'h22;
Memory[10872] = 8'hB3;
Memory[10879] = 8'h00;
Memory[10878] = 8'h02;
Memory[10877] = 8'h84;
Memory[10876] = 8'h63;
Memory[10883] = 8'h09;
Memory[10882] = 8'hD0;
Memory[10881] = 8'h50;
Memory[10880] = 8'h6F;
Memory[10887] = 8'h49;
Memory[10886] = 8'h8C;
Memory[10885] = 8'hA2;
Memory[10884] = 8'h03;
Memory[10891] = 8'h00;
Memory[10890] = 8'h32;
Memory[10889] = 8'h22;
Memory[10888] = 8'hB3;
Memory[10895] = 8'h00;
Memory[10894] = 8'h02;
Memory[10893] = 8'h84;
Memory[10892] = 8'h63;
Memory[10899] = 8'h09;
Memory[10898] = 8'h10;
Memory[10897] = 8'h50;
Memory[10896] = 8'h6F;
Memory[10903] = 8'h49;
Memory[10902] = 8'h4C;
Memory[10901] = 8'hA2;
Memory[10900] = 8'h03;
Memory[10907] = 8'h00;
Memory[10906] = 8'h32;
Memory[10905] = 8'h22;
Memory[10904] = 8'hB3;
Memory[10911] = 8'h00;
Memory[10910] = 8'h02;
Memory[10909] = 8'h84;
Memory[10908] = 8'h63;
Memory[10915] = 8'h08;
Memory[10914] = 8'h50;
Memory[10913] = 8'h50;
Memory[10912] = 8'h6F;
Memory[10919] = 8'h49;
Memory[10918] = 8'h0C;
Memory[10917] = 8'hA2;
Memory[10916] = 8'h03;
Memory[10923] = 8'h00;
Memory[10922] = 8'h32;
Memory[10921] = 8'h22;
Memory[10920] = 8'hB3;
Memory[10927] = 8'h00;
Memory[10926] = 8'h02;
Memory[10925] = 8'h84;
Memory[10924] = 8'h63;
Memory[10931] = 8'h07;
Memory[10930] = 8'h90;
Memory[10929] = 8'h50;
Memory[10928] = 8'h6F;
Memory[10935] = 8'h48;
Memory[10934] = 8'hCC;
Memory[10933] = 8'hA2;
Memory[10932] = 8'h03;
Memory[10939] = 8'h00;
Memory[10938] = 8'h32;
Memory[10937] = 8'h22;
Memory[10936] = 8'hB3;
Memory[10943] = 8'h00;
Memory[10942] = 8'h02;
Memory[10941] = 8'h84;
Memory[10940] = 8'h63;
Memory[10947] = 8'h06;
Memory[10946] = 8'hD0;
Memory[10945] = 8'h50;
Memory[10944] = 8'h6F;
Memory[10951] = 8'h48;
Memory[10950] = 8'h8C;
Memory[10949] = 8'hA2;
Memory[10948] = 8'h03;
Memory[10955] = 8'h00;
Memory[10954] = 8'h32;
Memory[10953] = 8'h22;
Memory[10952] = 8'hB3;
Memory[10959] = 8'h00;
Memory[10958] = 8'h02;
Memory[10957] = 8'h84;
Memory[10956] = 8'h63;
Memory[10963] = 8'h06;
Memory[10962] = 8'h10;
Memory[10961] = 8'h50;
Memory[10960] = 8'h6F;
Memory[10967] = 8'h48;
Memory[10966] = 8'h4C;
Memory[10965] = 8'hA2;
Memory[10964] = 8'h03;
Memory[10971] = 8'h00;
Memory[10970] = 8'h32;
Memory[10969] = 8'h22;
Memory[10968] = 8'hB3;
Memory[10975] = 8'h00;
Memory[10974] = 8'h02;
Memory[10973] = 8'h84;
Memory[10972] = 8'h63;
Memory[10979] = 8'h05;
Memory[10978] = 8'h50;
Memory[10977] = 8'h50;
Memory[10976] = 8'h6F;
Memory[10983] = 8'h48;
Memory[10982] = 8'h0C;
Memory[10981] = 8'hA2;
Memory[10980] = 8'h03;
Memory[10987] = 8'h00;
Memory[10986] = 8'h32;
Memory[10985] = 8'h22;
Memory[10984] = 8'hB3;
Memory[10991] = 8'h00;
Memory[10990] = 8'h02;
Memory[10989] = 8'h84;
Memory[10988] = 8'h63;
Memory[10995] = 8'h04;
Memory[10994] = 8'h90;
Memory[10993] = 8'h50;
Memory[10992] = 8'h6F;
Memory[10999] = 8'h47;
Memory[10998] = 8'hCC;
Memory[10997] = 8'hA2;
Memory[10996] = 8'h03;
Memory[11003] = 8'h00;
Memory[11002] = 8'h32;
Memory[11001] = 8'h22;
Memory[11000] = 8'hB3;
Memory[11007] = 8'h00;
Memory[11006] = 8'h02;
Memory[11005] = 8'h84;
Memory[11004] = 8'h63;
Memory[11011] = 8'h03;
Memory[11010] = 8'hD0;
Memory[11009] = 8'h50;
Memory[11008] = 8'h6F;
Memory[11015] = 8'h47;
Memory[11014] = 8'h8C;
Memory[11013] = 8'hA2;
Memory[11012] = 8'h03;
Memory[11019] = 8'h00;
Memory[11018] = 8'h32;
Memory[11017] = 8'h22;
Memory[11016] = 8'hB3;
Memory[11023] = 8'h00;
Memory[11022] = 8'h02;
Memory[11021] = 8'h84;
Memory[11020] = 8'h63;
Memory[11027] = 8'h03;
Memory[11026] = 8'h10;
Memory[11025] = 8'h50;
Memory[11024] = 8'h6F;
Memory[11031] = 8'h47;
Memory[11030] = 8'h4C;
Memory[11029] = 8'hA2;
Memory[11028] = 8'h03;
Memory[11035] = 8'h00;
Memory[11034] = 8'h32;
Memory[11033] = 8'h22;
Memory[11032] = 8'hB3;
Memory[11039] = 8'h00;
Memory[11038] = 8'h02;
Memory[11037] = 8'h84;
Memory[11036] = 8'h63;
Memory[11043] = 8'h02;
Memory[11042] = 8'h50;
Memory[11041] = 8'h50;
Memory[11040] = 8'h6F;
Memory[11047] = 8'h47;
Memory[11046] = 8'h0C;
Memory[11045] = 8'hA2;
Memory[11044] = 8'h03;
Memory[11051] = 8'h00;
Memory[11050] = 8'h32;
Memory[11049] = 8'h22;
Memory[11048] = 8'hB3;
Memory[11055] = 8'h00;
Memory[11054] = 8'h02;
Memory[11053] = 8'h84;
Memory[11052] = 8'h63;
Memory[11059] = 8'h01;
Memory[11058] = 8'h90;
Memory[11057] = 8'h50;
Memory[11056] = 8'h6F;
Memory[11063] = 8'h46;
Memory[11062] = 8'hCC;
Memory[11061] = 8'hA2;
Memory[11060] = 8'h03;
Memory[11067] = 8'h00;
Memory[11066] = 8'h32;
Memory[11065] = 8'h22;
Memory[11064] = 8'hB3;
Memory[11071] = 8'h00;
Memory[11070] = 8'h02;
Memory[11069] = 8'h84;
Memory[11068] = 8'h63;
Memory[11075] = 8'h00;
Memory[11074] = 8'hD0;
Memory[11073] = 8'h50;
Memory[11072] = 8'h6F;
Memory[11079] = 8'h46;
Memory[11078] = 8'h8C;
Memory[11077] = 8'hA2;
Memory[11076] = 8'h03;
Memory[11083] = 8'h00;
Memory[11082] = 8'h32;
Memory[11081] = 8'h22;
Memory[11080] = 8'hB3;
Memory[11087] = 8'h00;
Memory[11086] = 8'h02;
Memory[11085] = 8'h84;
Memory[11084] = 8'h63;
Memory[11091] = 8'h00;
Memory[11090] = 8'h10;
Memory[11089] = 8'h50;
Memory[11088] = 8'h6F;
Memory[11095] = 8'h46;
Memory[11094] = 8'h4C;
Memory[11093] = 8'hA2;
Memory[11092] = 8'h03;
Memory[11099] = 8'h00;
Memory[11098] = 8'h32;
Memory[11097] = 8'h22;
Memory[11096] = 8'hB3;
Memory[11103] = 8'h00;
Memory[11102] = 8'h02;
Memory[11101] = 8'h84;
Memory[11100] = 8'h63;
Memory[11107] = 8'h7F;
Memory[11106] = 8'h40;
Memory[11105] = 8'h50;
Memory[11104] = 8'h6F;
Memory[11111] = 8'h46;
Memory[11110] = 8'h0C;
Memory[11109] = 8'hA2;
Memory[11108] = 8'h03;
Memory[11115] = 8'h00;
Memory[11114] = 8'h32;
Memory[11113] = 8'h22;
Memory[11112] = 8'hB3;
Memory[11119] = 8'h00;
Memory[11118] = 8'h02;
Memory[11117] = 8'h84;
Memory[11116] = 8'h63;
Memory[11123] = 8'h7E;
Memory[11122] = 8'h80;
Memory[11121] = 8'h50;
Memory[11120] = 8'h6F;
Memory[11127] = 8'h45;
Memory[11126] = 8'hCC;
Memory[11125] = 8'hA2;
Memory[11124] = 8'h03;
Memory[11131] = 8'h00;
Memory[11130] = 8'h32;
Memory[11129] = 8'h22;
Memory[11128] = 8'hB3;
Memory[11135] = 8'h00;
Memory[11134] = 8'h02;
Memory[11133] = 8'h84;
Memory[11132] = 8'h63;
Memory[11139] = 8'h7D;
Memory[11138] = 8'hC0;
Memory[11137] = 8'h50;
Memory[11136] = 8'h6F;
Memory[11143] = 8'h45;
Memory[11142] = 8'h8C;
Memory[11141] = 8'hA2;
Memory[11140] = 8'h03;
Memory[11147] = 8'h00;
Memory[11146] = 8'h32;
Memory[11145] = 8'h22;
Memory[11144] = 8'hB3;
Memory[11151] = 8'h00;
Memory[11150] = 8'h02;
Memory[11149] = 8'h84;
Memory[11148] = 8'h63;
Memory[11155] = 8'h7D;
Memory[11154] = 8'h00;
Memory[11153] = 8'h50;
Memory[11152] = 8'h6F;
Memory[11159] = 8'h45;
Memory[11158] = 8'h4C;
Memory[11157] = 8'hA2;
Memory[11156] = 8'h03;
Memory[11163] = 8'h00;
Memory[11162] = 8'h32;
Memory[11161] = 8'h22;
Memory[11160] = 8'hB3;
Memory[11167] = 8'h00;
Memory[11166] = 8'h02;
Memory[11165] = 8'h84;
Memory[11164] = 8'h63;
Memory[11171] = 8'h7C;
Memory[11170] = 8'h40;
Memory[11169] = 8'h50;
Memory[11168] = 8'h6F;
Memory[11175] = 8'h45;
Memory[11174] = 8'h0C;
Memory[11173] = 8'hA2;
Memory[11172] = 8'h03;
Memory[11179] = 8'h00;
Memory[11178] = 8'h32;
Memory[11177] = 8'h22;
Memory[11176] = 8'hB3;
Memory[11183] = 8'h00;
Memory[11182] = 8'h02;
Memory[11181] = 8'h84;
Memory[11180] = 8'h63;
Memory[11187] = 8'h7B;
Memory[11186] = 8'h80;
Memory[11185] = 8'h50;
Memory[11184] = 8'h6F;
Memory[11191] = 8'h44;
Memory[11190] = 8'hCC;
Memory[11189] = 8'hA2;
Memory[11188] = 8'h03;
Memory[11195] = 8'h00;
Memory[11194] = 8'h32;
Memory[11193] = 8'h22;
Memory[11192] = 8'hB3;
Memory[11199] = 8'h00;
Memory[11198] = 8'h02;
Memory[11197] = 8'h84;
Memory[11196] = 8'h63;
Memory[11203] = 8'h7A;
Memory[11202] = 8'hC0;
Memory[11201] = 8'h50;
Memory[11200] = 8'h6F;
Memory[11207] = 8'h44;
Memory[11206] = 8'h8C;
Memory[11205] = 8'hA2;
Memory[11204] = 8'h03;
Memory[11211] = 8'h00;
Memory[11210] = 8'h32;
Memory[11209] = 8'h22;
Memory[11208] = 8'hB3;
Memory[11215] = 8'h00;
Memory[11214] = 8'h02;
Memory[11213] = 8'h84;
Memory[11212] = 8'h63;
Memory[11219] = 8'h7A;
Memory[11218] = 8'h00;
Memory[11217] = 8'h50;
Memory[11216] = 8'h6F;
Memory[11223] = 8'h44;
Memory[11222] = 8'h4C;
Memory[11221] = 8'hA2;
Memory[11220] = 8'h03;
Memory[11227] = 8'h00;
Memory[11226] = 8'h32;
Memory[11225] = 8'h22;
Memory[11224] = 8'hB3;
Memory[11231] = 8'h00;
Memory[11230] = 8'h02;
Memory[11229] = 8'h84;
Memory[11228] = 8'h63;
Memory[11235] = 8'h79;
Memory[11234] = 8'h40;
Memory[11233] = 8'h50;
Memory[11232] = 8'h6F;
Memory[11239] = 8'h44;
Memory[11238] = 8'h0C;
Memory[11237] = 8'hA2;
Memory[11236] = 8'h03;
Memory[11243] = 8'h00;
Memory[11242] = 8'h32;
Memory[11241] = 8'h22;
Memory[11240] = 8'hB3;
Memory[11247] = 8'h00;
Memory[11246] = 8'h02;
Memory[11245] = 8'h84;
Memory[11244] = 8'h63;
Memory[11251] = 8'h78;
Memory[11250] = 8'h80;
Memory[11249] = 8'h50;
Memory[11248] = 8'h6F;
Memory[11255] = 8'h43;
Memory[11254] = 8'hCC;
Memory[11253] = 8'hA2;
Memory[11252] = 8'h03;
Memory[11259] = 8'h00;
Memory[11258] = 8'h32;
Memory[11257] = 8'h22;
Memory[11256] = 8'hB3;
Memory[11263] = 8'h00;
Memory[11262] = 8'h02;
Memory[11261] = 8'h84;
Memory[11260] = 8'h63;
Memory[11267] = 8'h77;
Memory[11266] = 8'hC0;
Memory[11265] = 8'h50;
Memory[11264] = 8'h6F;
Memory[11271] = 8'h43;
Memory[11270] = 8'h8C;
Memory[11269] = 8'hA2;
Memory[11268] = 8'h03;
Memory[11275] = 8'h00;
Memory[11274] = 8'h32;
Memory[11273] = 8'h22;
Memory[11272] = 8'hB3;
Memory[11279] = 8'h00;
Memory[11278] = 8'h02;
Memory[11277] = 8'h84;
Memory[11276] = 8'h63;
Memory[11283] = 8'h77;
Memory[11282] = 8'h00;
Memory[11281] = 8'h50;
Memory[11280] = 8'h6F;
Memory[11287] = 8'h43;
Memory[11286] = 8'h4C;
Memory[11285] = 8'hA2;
Memory[11284] = 8'h03;
Memory[11291] = 8'h00;
Memory[11290] = 8'h32;
Memory[11289] = 8'h22;
Memory[11288] = 8'hB3;
Memory[11295] = 8'h00;
Memory[11294] = 8'h02;
Memory[11293] = 8'h84;
Memory[11292] = 8'h63;
Memory[11299] = 8'h76;
Memory[11298] = 8'h40;
Memory[11297] = 8'h50;
Memory[11296] = 8'h6F;
Memory[11303] = 8'h43;
Memory[11302] = 8'h0C;
Memory[11301] = 8'hA2;
Memory[11300] = 8'h03;
Memory[11307] = 8'h00;
Memory[11306] = 8'h32;
Memory[11305] = 8'h22;
Memory[11304] = 8'hB3;
Memory[11311] = 8'h00;
Memory[11310] = 8'h02;
Memory[11309] = 8'h84;
Memory[11308] = 8'h63;
Memory[11315] = 8'h75;
Memory[11314] = 8'h80;
Memory[11313] = 8'h50;
Memory[11312] = 8'h6F;
Memory[11319] = 8'h42;
Memory[11318] = 8'hCC;
Memory[11317] = 8'hA2;
Memory[11316] = 8'h03;
Memory[11323] = 8'h00;
Memory[11322] = 8'h32;
Memory[11321] = 8'h22;
Memory[11320] = 8'hB3;
Memory[11327] = 8'h00;
Memory[11326] = 8'h02;
Memory[11325] = 8'h84;
Memory[11324] = 8'h63;
Memory[11331] = 8'h74;
Memory[11330] = 8'hC0;
Memory[11329] = 8'h50;
Memory[11328] = 8'h6F;
Memory[11335] = 8'h42;
Memory[11334] = 8'h8C;
Memory[11333] = 8'hA2;
Memory[11332] = 8'h03;
Memory[11339] = 8'h00;
Memory[11338] = 8'h32;
Memory[11337] = 8'h22;
Memory[11336] = 8'hB3;
Memory[11343] = 8'h00;
Memory[11342] = 8'h02;
Memory[11341] = 8'h84;
Memory[11340] = 8'h63;
Memory[11347] = 8'h74;
Memory[11346] = 8'h00;
Memory[11345] = 8'h50;
Memory[11344] = 8'h6F;
Memory[11351] = 8'h42;
Memory[11350] = 8'h4C;
Memory[11349] = 8'hA2;
Memory[11348] = 8'h03;
Memory[11355] = 8'h00;
Memory[11354] = 8'h32;
Memory[11353] = 8'h22;
Memory[11352] = 8'hB3;
Memory[11359] = 8'h00;
Memory[11358] = 8'h02;
Memory[11357] = 8'h84;
Memory[11356] = 8'h63;
Memory[11363] = 8'h73;
Memory[11362] = 8'h40;
Memory[11361] = 8'h50;
Memory[11360] = 8'h6F;
Memory[11367] = 8'h42;
Memory[11366] = 8'h0C;
Memory[11365] = 8'hA2;
Memory[11364] = 8'h03;
Memory[11371] = 8'h00;
Memory[11370] = 8'h32;
Memory[11369] = 8'h22;
Memory[11368] = 8'hB3;
Memory[11375] = 8'h00;
Memory[11374] = 8'h02;
Memory[11373] = 8'h84;
Memory[11372] = 8'h63;
Memory[11379] = 8'h72;
Memory[11378] = 8'h80;
Memory[11377] = 8'h50;
Memory[11376] = 8'h6F;
Memory[11383] = 8'h41;
Memory[11382] = 8'hCC;
Memory[11381] = 8'hA2;
Memory[11380] = 8'h03;
Memory[11387] = 8'h00;
Memory[11386] = 8'h32;
Memory[11385] = 8'h22;
Memory[11384] = 8'hB3;
Memory[11391] = 8'h00;
Memory[11390] = 8'h02;
Memory[11389] = 8'h84;
Memory[11388] = 8'h63;
Memory[11395] = 8'h71;
Memory[11394] = 8'hC0;
Memory[11393] = 8'h50;
Memory[11392] = 8'h6F;
Memory[11399] = 8'h41;
Memory[11398] = 8'h8C;
Memory[11397] = 8'hA2;
Memory[11396] = 8'h03;
Memory[11403] = 8'h00;
Memory[11402] = 8'h32;
Memory[11401] = 8'h22;
Memory[11400] = 8'hB3;
Memory[11407] = 8'h00;
Memory[11406] = 8'h02;
Memory[11405] = 8'h84;
Memory[11404] = 8'h63;
Memory[11411] = 8'h71;
Memory[11410] = 8'h00;
Memory[11409] = 8'h50;
Memory[11408] = 8'h6F;
Memory[11415] = 8'h41;
Memory[11414] = 8'h4C;
Memory[11413] = 8'hA2;
Memory[11412] = 8'h03;
Memory[11419] = 8'h00;
Memory[11418] = 8'h32;
Memory[11417] = 8'h22;
Memory[11416] = 8'hB3;
Memory[11423] = 8'h00;
Memory[11422] = 8'h02;
Memory[11421] = 8'h84;
Memory[11420] = 8'h63;
Memory[11427] = 8'h70;
Memory[11426] = 8'h40;
Memory[11425] = 8'h50;
Memory[11424] = 8'h6F;
Memory[11431] = 8'h41;
Memory[11430] = 8'h0C;
Memory[11429] = 8'hA2;
Memory[11428] = 8'h03;
Memory[11435] = 8'h00;
Memory[11434] = 8'h32;
Memory[11433] = 8'h22;
Memory[11432] = 8'hB3;
Memory[11439] = 8'h00;
Memory[11438] = 8'h02;
Memory[11437] = 8'h84;
Memory[11436] = 8'h63;
Memory[11443] = 8'h6F;
Memory[11442] = 8'h80;
Memory[11441] = 8'h50;
Memory[11440] = 8'h6F;
Memory[11447] = 8'h40;
Memory[11446] = 8'hCC;
Memory[11445] = 8'hA2;
Memory[11444] = 8'h03;
Memory[11451] = 8'h00;
Memory[11450] = 8'h32;
Memory[11449] = 8'h22;
Memory[11448] = 8'hB3;
Memory[11455] = 8'h00;
Memory[11454] = 8'h02;
Memory[11453] = 8'h84;
Memory[11452] = 8'h63;
Memory[11459] = 8'h6E;
Memory[11458] = 8'hC0;
Memory[11457] = 8'h50;
Memory[11456] = 8'h6F;
Memory[11463] = 8'h40;
Memory[11462] = 8'h8C;
Memory[11461] = 8'hA2;
Memory[11460] = 8'h03;
Memory[11467] = 8'h00;
Memory[11466] = 8'h32;
Memory[11465] = 8'h22;
Memory[11464] = 8'hB3;
Memory[11471] = 8'h00;
Memory[11470] = 8'h02;
Memory[11469] = 8'h84;
Memory[11468] = 8'h63;
Memory[11475] = 8'h6E;
Memory[11474] = 8'h00;
Memory[11473] = 8'h50;
Memory[11472] = 8'h6F;
Memory[11479] = 8'h40;
Memory[11478] = 8'h4C;
Memory[11477] = 8'hA2;
Memory[11476] = 8'h03;
Memory[11483] = 8'h00;
Memory[11482] = 8'h32;
Memory[11481] = 8'h22;
Memory[11480] = 8'hB3;
Memory[11487] = 8'h00;
Memory[11486] = 8'h02;
Memory[11485] = 8'h84;
Memory[11484] = 8'h63;
Memory[11491] = 8'h6D;
Memory[11490] = 8'h40;
Memory[11489] = 8'h50;
Memory[11488] = 8'h6F;
Memory[11495] = 8'h40;
Memory[11494] = 8'h0C;
Memory[11493] = 8'hA2;
Memory[11492] = 8'h03;
Memory[11499] = 8'h00;
Memory[11498] = 8'h32;
Memory[11497] = 8'h22;
Memory[11496] = 8'hB3;
Memory[11503] = 8'h00;
Memory[11502] = 8'h02;
Memory[11501] = 8'h84;
Memory[11500] = 8'h63;
Memory[11507] = 8'h6C;
Memory[11506] = 8'h80;
Memory[11505] = 8'h50;
Memory[11504] = 8'h6F;
Memory[11511] = 8'h3F;
Memory[11510] = 8'hCC;
Memory[11509] = 8'hA2;
Memory[11508] = 8'h03;
Memory[11515] = 8'h00;
Memory[11514] = 8'h32;
Memory[11513] = 8'h22;
Memory[11512] = 8'hB3;
Memory[11519] = 8'h00;
Memory[11518] = 8'h02;
Memory[11517] = 8'h84;
Memory[11516] = 8'h63;
Memory[11523] = 8'h6B;
Memory[11522] = 8'hC0;
Memory[11521] = 8'h50;
Memory[11520] = 8'h6F;
Memory[11527] = 8'h3F;
Memory[11526] = 8'h8C;
Memory[11525] = 8'hA2;
Memory[11524] = 8'h03;
Memory[11531] = 8'h00;
Memory[11530] = 8'h32;
Memory[11529] = 8'h22;
Memory[11528] = 8'hB3;
Memory[11535] = 8'h00;
Memory[11534] = 8'h02;
Memory[11533] = 8'h84;
Memory[11532] = 8'h63;
Memory[11539] = 8'h6B;
Memory[11538] = 8'h00;
Memory[11537] = 8'h50;
Memory[11536] = 8'h6F;
Memory[11543] = 8'h3F;
Memory[11542] = 8'h4C;
Memory[11541] = 8'hA2;
Memory[11540] = 8'h03;
Memory[11547] = 8'h00;
Memory[11546] = 8'h32;
Memory[11545] = 8'h22;
Memory[11544] = 8'hB3;
Memory[11551] = 8'h00;
Memory[11550] = 8'h02;
Memory[11549] = 8'h84;
Memory[11548] = 8'h63;
Memory[11555] = 8'h6A;
Memory[11554] = 8'h40;
Memory[11553] = 8'h50;
Memory[11552] = 8'h6F;
Memory[11559] = 8'h3F;
Memory[11558] = 8'h0C;
Memory[11557] = 8'hA2;
Memory[11556] = 8'h03;
Memory[11563] = 8'h00;
Memory[11562] = 8'h32;
Memory[11561] = 8'h22;
Memory[11560] = 8'hB3;
Memory[11567] = 8'h00;
Memory[11566] = 8'h02;
Memory[11565] = 8'h84;
Memory[11564] = 8'h63;
Memory[11571] = 8'h69;
Memory[11570] = 8'h80;
Memory[11569] = 8'h50;
Memory[11568] = 8'h6F;
Memory[11575] = 8'h3E;
Memory[11574] = 8'hCC;
Memory[11573] = 8'hA2;
Memory[11572] = 8'h03;
Memory[11579] = 8'h00;
Memory[11578] = 8'h32;
Memory[11577] = 8'h22;
Memory[11576] = 8'hB3;
Memory[11583] = 8'h00;
Memory[11582] = 8'h02;
Memory[11581] = 8'h84;
Memory[11580] = 8'h63;
Memory[11587] = 8'h68;
Memory[11586] = 8'hC0;
Memory[11585] = 8'h50;
Memory[11584] = 8'h6F;
Memory[11591] = 8'h3E;
Memory[11590] = 8'h8C;
Memory[11589] = 8'hA2;
Memory[11588] = 8'h03;
Memory[11595] = 8'h00;
Memory[11594] = 8'h32;
Memory[11593] = 8'h22;
Memory[11592] = 8'hB3;
Memory[11599] = 8'h00;
Memory[11598] = 8'h02;
Memory[11597] = 8'h84;
Memory[11596] = 8'h63;
Memory[11603] = 8'h68;
Memory[11602] = 8'h00;
Memory[11601] = 8'h50;
Memory[11600] = 8'h6F;
Memory[11607] = 8'h3E;
Memory[11606] = 8'h4C;
Memory[11605] = 8'hA2;
Memory[11604] = 8'h03;
Memory[11611] = 8'h00;
Memory[11610] = 8'h32;
Memory[11609] = 8'h22;
Memory[11608] = 8'hB3;
Memory[11615] = 8'h00;
Memory[11614] = 8'h02;
Memory[11613] = 8'h84;
Memory[11612] = 8'h63;
Memory[11619] = 8'h67;
Memory[11618] = 8'h40;
Memory[11617] = 8'h50;
Memory[11616] = 8'h6F;
Memory[11623] = 8'h3E;
Memory[11622] = 8'h0C;
Memory[11621] = 8'hA2;
Memory[11620] = 8'h03;
Memory[11627] = 8'h00;
Memory[11626] = 8'h32;
Memory[11625] = 8'h22;
Memory[11624] = 8'hB3;
Memory[11631] = 8'h00;
Memory[11630] = 8'h02;
Memory[11629] = 8'h84;
Memory[11628] = 8'h63;
Memory[11635] = 8'h66;
Memory[11634] = 8'h80;
Memory[11633] = 8'h50;
Memory[11632] = 8'h6F;
Memory[11639] = 8'h3D;
Memory[11638] = 8'hCC;
Memory[11637] = 8'hA2;
Memory[11636] = 8'h03;
Memory[11643] = 8'h00;
Memory[11642] = 8'h32;
Memory[11641] = 8'h22;
Memory[11640] = 8'hB3;
Memory[11647] = 8'h00;
Memory[11646] = 8'h02;
Memory[11645] = 8'h84;
Memory[11644] = 8'h63;
Memory[11651] = 8'h65;
Memory[11650] = 8'hC0;
Memory[11649] = 8'h50;
Memory[11648] = 8'h6F;
Memory[11655] = 8'h3D;
Memory[11654] = 8'h8C;
Memory[11653] = 8'hA2;
Memory[11652] = 8'h03;
Memory[11659] = 8'h00;
Memory[11658] = 8'h32;
Memory[11657] = 8'h22;
Memory[11656] = 8'hB3;
Memory[11663] = 8'h00;
Memory[11662] = 8'h02;
Memory[11661] = 8'h84;
Memory[11660] = 8'h63;
Memory[11667] = 8'h65;
Memory[11666] = 8'h00;
Memory[11665] = 8'h50;
Memory[11664] = 8'h6F;
Memory[11671] = 8'h3D;
Memory[11670] = 8'h4C;
Memory[11669] = 8'hA2;
Memory[11668] = 8'h03;
Memory[11675] = 8'h00;
Memory[11674] = 8'h32;
Memory[11673] = 8'h22;
Memory[11672] = 8'hB3;
Memory[11679] = 8'h00;
Memory[11678] = 8'h02;
Memory[11677] = 8'h84;
Memory[11676] = 8'h63;
Memory[11683] = 8'h64;
Memory[11682] = 8'h40;
Memory[11681] = 8'h50;
Memory[11680] = 8'h6F;
Memory[11687] = 8'h3D;
Memory[11686] = 8'h0C;
Memory[11685] = 8'hA2;
Memory[11684] = 8'h03;
Memory[11691] = 8'h00;
Memory[11690] = 8'h32;
Memory[11689] = 8'h22;
Memory[11688] = 8'hB3;
Memory[11695] = 8'h00;
Memory[11694] = 8'h02;
Memory[11693] = 8'h84;
Memory[11692] = 8'h63;
Memory[11699] = 8'h63;
Memory[11698] = 8'h80;
Memory[11697] = 8'h50;
Memory[11696] = 8'h6F;
Memory[11703] = 8'h3C;
Memory[11702] = 8'hCC;
Memory[11701] = 8'hA2;
Memory[11700] = 8'h03;
Memory[11707] = 8'h00;
Memory[11706] = 8'h32;
Memory[11705] = 8'h22;
Memory[11704] = 8'hB3;
Memory[11711] = 8'h00;
Memory[11710] = 8'h02;
Memory[11709] = 8'h84;
Memory[11708] = 8'h63;
Memory[11715] = 8'h62;
Memory[11714] = 8'hC0;
Memory[11713] = 8'h50;
Memory[11712] = 8'h6F;
Memory[11719] = 8'h3C;
Memory[11718] = 8'h8C;
Memory[11717] = 8'hA2;
Memory[11716] = 8'h03;
Memory[11723] = 8'h00;
Memory[11722] = 8'h32;
Memory[11721] = 8'h22;
Memory[11720] = 8'hB3;
Memory[11727] = 8'h00;
Memory[11726] = 8'h02;
Memory[11725] = 8'h84;
Memory[11724] = 8'h63;
Memory[11731] = 8'h62;
Memory[11730] = 8'h00;
Memory[11729] = 8'h50;
Memory[11728] = 8'h6F;
Memory[11735] = 8'h3C;
Memory[11734] = 8'h4C;
Memory[11733] = 8'hA2;
Memory[11732] = 8'h03;
Memory[11739] = 8'h00;
Memory[11738] = 8'h32;
Memory[11737] = 8'h22;
Memory[11736] = 8'hB3;
Memory[11743] = 8'h00;
Memory[11742] = 8'h02;
Memory[11741] = 8'h84;
Memory[11740] = 8'h63;
Memory[11747] = 8'h61;
Memory[11746] = 8'h40;
Memory[11745] = 8'h50;
Memory[11744] = 8'h6F;
Memory[11751] = 8'h3C;
Memory[11750] = 8'h0C;
Memory[11749] = 8'hA2;
Memory[11748] = 8'h03;
Memory[11755] = 8'h00;
Memory[11754] = 8'h32;
Memory[11753] = 8'h22;
Memory[11752] = 8'hB3;
Memory[11759] = 8'h00;
Memory[11758] = 8'h02;
Memory[11757] = 8'h84;
Memory[11756] = 8'h63;
Memory[11763] = 8'h60;
Memory[11762] = 8'h80;
Memory[11761] = 8'h50;
Memory[11760] = 8'h6F;
Memory[11767] = 8'h3B;
Memory[11766] = 8'hCC;
Memory[11765] = 8'hA2;
Memory[11764] = 8'h03;
Memory[11771] = 8'h00;
Memory[11770] = 8'h32;
Memory[11769] = 8'h22;
Memory[11768] = 8'hB3;
Memory[11775] = 8'h00;
Memory[11774] = 8'h02;
Memory[11773] = 8'h84;
Memory[11772] = 8'h63;
Memory[11779] = 8'h5F;
Memory[11778] = 8'hC0;
Memory[11777] = 8'h50;
Memory[11776] = 8'h6F;
Memory[11783] = 8'h3B;
Memory[11782] = 8'h8C;
Memory[11781] = 8'hA2;
Memory[11780] = 8'h03;
Memory[11787] = 8'h00;
Memory[11786] = 8'h32;
Memory[11785] = 8'h22;
Memory[11784] = 8'hB3;
Memory[11791] = 8'h00;
Memory[11790] = 8'h02;
Memory[11789] = 8'h84;
Memory[11788] = 8'h63;
Memory[11795] = 8'h5F;
Memory[11794] = 8'h00;
Memory[11793] = 8'h50;
Memory[11792] = 8'h6F;
Memory[11799] = 8'h3B;
Memory[11798] = 8'h4C;
Memory[11797] = 8'hA2;
Memory[11796] = 8'h03;
Memory[11803] = 8'h00;
Memory[11802] = 8'h32;
Memory[11801] = 8'h22;
Memory[11800] = 8'hB3;
Memory[11807] = 8'h00;
Memory[11806] = 8'h02;
Memory[11805] = 8'h84;
Memory[11804] = 8'h63;
Memory[11811] = 8'h5E;
Memory[11810] = 8'h40;
Memory[11809] = 8'h50;
Memory[11808] = 8'h6F;
Memory[11815] = 8'h3B;
Memory[11814] = 8'h0C;
Memory[11813] = 8'hA2;
Memory[11812] = 8'h03;
Memory[11819] = 8'h00;
Memory[11818] = 8'h32;
Memory[11817] = 8'h22;
Memory[11816] = 8'hB3;
Memory[11823] = 8'h00;
Memory[11822] = 8'h02;
Memory[11821] = 8'h84;
Memory[11820] = 8'h63;
Memory[11827] = 8'h5D;
Memory[11826] = 8'h80;
Memory[11825] = 8'h50;
Memory[11824] = 8'h6F;
Memory[11831] = 8'h3A;
Memory[11830] = 8'hCC;
Memory[11829] = 8'hA2;
Memory[11828] = 8'h03;
Memory[11835] = 8'h00;
Memory[11834] = 8'h32;
Memory[11833] = 8'h22;
Memory[11832] = 8'hB3;
Memory[11839] = 8'h00;
Memory[11838] = 8'h02;
Memory[11837] = 8'h84;
Memory[11836] = 8'h63;
Memory[11843] = 8'h5C;
Memory[11842] = 8'hC0;
Memory[11841] = 8'h50;
Memory[11840] = 8'h6F;
Memory[11847] = 8'h3A;
Memory[11846] = 8'h8C;
Memory[11845] = 8'hA2;
Memory[11844] = 8'h03;
Memory[11851] = 8'h00;
Memory[11850] = 8'h32;
Memory[11849] = 8'h22;
Memory[11848] = 8'hB3;
Memory[11855] = 8'h00;
Memory[11854] = 8'h02;
Memory[11853] = 8'h84;
Memory[11852] = 8'h63;
Memory[11859] = 8'h5C;
Memory[11858] = 8'h00;
Memory[11857] = 8'h50;
Memory[11856] = 8'h6F;
Memory[11863] = 8'h3A;
Memory[11862] = 8'h4C;
Memory[11861] = 8'hA2;
Memory[11860] = 8'h03;
Memory[11867] = 8'h00;
Memory[11866] = 8'h32;
Memory[11865] = 8'h22;
Memory[11864] = 8'hB3;
Memory[11871] = 8'h00;
Memory[11870] = 8'h02;
Memory[11869] = 8'h84;
Memory[11868] = 8'h63;
Memory[11875] = 8'h5B;
Memory[11874] = 8'h40;
Memory[11873] = 8'h50;
Memory[11872] = 8'h6F;
Memory[11879] = 8'h3A;
Memory[11878] = 8'h0C;
Memory[11877] = 8'hA2;
Memory[11876] = 8'h03;
Memory[11883] = 8'h00;
Memory[11882] = 8'h32;
Memory[11881] = 8'h22;
Memory[11880] = 8'hB3;
Memory[11887] = 8'h00;
Memory[11886] = 8'h02;
Memory[11885] = 8'h84;
Memory[11884] = 8'h63;
Memory[11891] = 8'h5A;
Memory[11890] = 8'h80;
Memory[11889] = 8'h50;
Memory[11888] = 8'h6F;
Memory[11895] = 8'h39;
Memory[11894] = 8'hCC;
Memory[11893] = 8'hA2;
Memory[11892] = 8'h03;
Memory[11899] = 8'h00;
Memory[11898] = 8'h32;
Memory[11897] = 8'h22;
Memory[11896] = 8'hB3;
Memory[11903] = 8'h00;
Memory[11902] = 8'h02;
Memory[11901] = 8'h84;
Memory[11900] = 8'h63;
Memory[11907] = 8'h59;
Memory[11906] = 8'hC0;
Memory[11905] = 8'h50;
Memory[11904] = 8'h6F;
Memory[11911] = 8'h39;
Memory[11910] = 8'h8C;
Memory[11909] = 8'hA2;
Memory[11908] = 8'h03;
Memory[11915] = 8'h00;
Memory[11914] = 8'h32;
Memory[11913] = 8'h22;
Memory[11912] = 8'hB3;
Memory[11919] = 8'h00;
Memory[11918] = 8'h02;
Memory[11917] = 8'h84;
Memory[11916] = 8'h63;
Memory[11923] = 8'h59;
Memory[11922] = 8'h00;
Memory[11921] = 8'h50;
Memory[11920] = 8'h6F;
Memory[11927] = 8'h39;
Memory[11926] = 8'h4C;
Memory[11925] = 8'hA2;
Memory[11924] = 8'h03;
Memory[11931] = 8'h00;
Memory[11930] = 8'h32;
Memory[11929] = 8'h22;
Memory[11928] = 8'hB3;
Memory[11935] = 8'h00;
Memory[11934] = 8'h02;
Memory[11933] = 8'h84;
Memory[11932] = 8'h63;
Memory[11939] = 8'h58;
Memory[11938] = 8'h40;
Memory[11937] = 8'h50;
Memory[11936] = 8'h6F;
Memory[11943] = 8'h39;
Memory[11942] = 8'h0C;
Memory[11941] = 8'hA2;
Memory[11940] = 8'h03;
Memory[11947] = 8'h00;
Memory[11946] = 8'h32;
Memory[11945] = 8'h22;
Memory[11944] = 8'hB3;
Memory[11951] = 8'h00;
Memory[11950] = 8'h02;
Memory[11949] = 8'h84;
Memory[11948] = 8'h63;
Memory[11955] = 8'h57;
Memory[11954] = 8'h80;
Memory[11953] = 8'h50;
Memory[11952] = 8'h6F;
Memory[11959] = 8'h38;
Memory[11958] = 8'hCC;
Memory[11957] = 8'hA2;
Memory[11956] = 8'h03;
Memory[11963] = 8'h00;
Memory[11962] = 8'h32;
Memory[11961] = 8'h22;
Memory[11960] = 8'hB3;
Memory[11967] = 8'h00;
Memory[11966] = 8'h02;
Memory[11965] = 8'h84;
Memory[11964] = 8'h63;
Memory[11971] = 8'h56;
Memory[11970] = 8'hC0;
Memory[11969] = 8'h50;
Memory[11968] = 8'h6F;
Memory[11975] = 8'h38;
Memory[11974] = 8'h8C;
Memory[11973] = 8'hA2;
Memory[11972] = 8'h03;
Memory[11979] = 8'h00;
Memory[11978] = 8'h32;
Memory[11977] = 8'h22;
Memory[11976] = 8'hB3;
Memory[11983] = 8'h00;
Memory[11982] = 8'h02;
Memory[11981] = 8'h84;
Memory[11980] = 8'h63;
Memory[11987] = 8'h56;
Memory[11986] = 8'h00;
Memory[11985] = 8'h50;
Memory[11984] = 8'h6F;
Memory[11991] = 8'h38;
Memory[11990] = 8'h4C;
Memory[11989] = 8'hA2;
Memory[11988] = 8'h03;
Memory[11995] = 8'h00;
Memory[11994] = 8'h32;
Memory[11993] = 8'h22;
Memory[11992] = 8'hB3;
Memory[11999] = 8'h00;
Memory[11998] = 8'h02;
Memory[11997] = 8'h84;
Memory[11996] = 8'h63;
Memory[12003] = 8'h55;
Memory[12002] = 8'h40;
Memory[12001] = 8'h50;
Memory[12000] = 8'h6F;
Memory[12007] = 8'h38;
Memory[12006] = 8'h0C;
Memory[12005] = 8'hA2;
Memory[12004] = 8'h03;
Memory[12011] = 8'h00;
Memory[12010] = 8'h32;
Memory[12009] = 8'h22;
Memory[12008] = 8'hB3;
Memory[12015] = 8'h00;
Memory[12014] = 8'h02;
Memory[12013] = 8'h84;
Memory[12012] = 8'h63;
Memory[12019] = 8'h54;
Memory[12018] = 8'h80;
Memory[12017] = 8'h50;
Memory[12016] = 8'h6F;
Memory[12023] = 8'h37;
Memory[12022] = 8'hCC;
Memory[12021] = 8'hA2;
Memory[12020] = 8'h03;
Memory[12027] = 8'h00;
Memory[12026] = 8'h32;
Memory[12025] = 8'h22;
Memory[12024] = 8'hB3;
Memory[12031] = 8'h00;
Memory[12030] = 8'h02;
Memory[12029] = 8'h84;
Memory[12028] = 8'h63;
Memory[12035] = 8'h53;
Memory[12034] = 8'hC0;
Memory[12033] = 8'h50;
Memory[12032] = 8'h6F;
Memory[12039] = 8'h37;
Memory[12038] = 8'h8C;
Memory[12037] = 8'hA2;
Memory[12036] = 8'h03;
Memory[12043] = 8'h00;
Memory[12042] = 8'h32;
Memory[12041] = 8'h22;
Memory[12040] = 8'hB3;
Memory[12047] = 8'h00;
Memory[12046] = 8'h02;
Memory[12045] = 8'h84;
Memory[12044] = 8'h63;
Memory[12051] = 8'h53;
Memory[12050] = 8'h00;
Memory[12049] = 8'h50;
Memory[12048] = 8'h6F;
Memory[12055] = 8'h37;
Memory[12054] = 8'h4C;
Memory[12053] = 8'hA2;
Memory[12052] = 8'h03;
Memory[12059] = 8'h00;
Memory[12058] = 8'h32;
Memory[12057] = 8'h22;
Memory[12056] = 8'hB3;
Memory[12063] = 8'h00;
Memory[12062] = 8'h02;
Memory[12061] = 8'h84;
Memory[12060] = 8'h63;
Memory[12067] = 8'h52;
Memory[12066] = 8'h40;
Memory[12065] = 8'h50;
Memory[12064] = 8'h6F;
Memory[12071] = 8'h37;
Memory[12070] = 8'h0C;
Memory[12069] = 8'hA2;
Memory[12068] = 8'h03;
Memory[12075] = 8'h00;
Memory[12074] = 8'h32;
Memory[12073] = 8'h22;
Memory[12072] = 8'hB3;
Memory[12079] = 8'h00;
Memory[12078] = 8'h02;
Memory[12077] = 8'h84;
Memory[12076] = 8'h63;
Memory[12083] = 8'h51;
Memory[12082] = 8'h80;
Memory[12081] = 8'h50;
Memory[12080] = 8'h6F;
Memory[12087] = 8'h36;
Memory[12086] = 8'hCC;
Memory[12085] = 8'hA2;
Memory[12084] = 8'h03;
Memory[12091] = 8'h00;
Memory[12090] = 8'h32;
Memory[12089] = 8'h22;
Memory[12088] = 8'hB3;
Memory[12095] = 8'h00;
Memory[12094] = 8'h02;
Memory[12093] = 8'h84;
Memory[12092] = 8'h63;
Memory[12099] = 8'h50;
Memory[12098] = 8'hC0;
Memory[12097] = 8'h50;
Memory[12096] = 8'h6F;
Memory[12103] = 8'h36;
Memory[12102] = 8'h8C;
Memory[12101] = 8'hA2;
Memory[12100] = 8'h03;
Memory[12107] = 8'h00;
Memory[12106] = 8'h32;
Memory[12105] = 8'h22;
Memory[12104] = 8'hB3;
Memory[12111] = 8'h00;
Memory[12110] = 8'h02;
Memory[12109] = 8'h84;
Memory[12108] = 8'h63;
Memory[12115] = 8'h50;
Memory[12114] = 8'h00;
Memory[12113] = 8'h50;
Memory[12112] = 8'h6F;
Memory[12119] = 8'h36;
Memory[12118] = 8'h4C;
Memory[12117] = 8'hA2;
Memory[12116] = 8'h03;
Memory[12123] = 8'h00;
Memory[12122] = 8'h32;
Memory[12121] = 8'h22;
Memory[12120] = 8'hB3;
Memory[12127] = 8'h00;
Memory[12126] = 8'h02;
Memory[12125] = 8'h84;
Memory[12124] = 8'h63;
Memory[12131] = 8'h4F;
Memory[12130] = 8'h40;
Memory[12129] = 8'h50;
Memory[12128] = 8'h6F;
Memory[12135] = 8'h36;
Memory[12134] = 8'h0C;
Memory[12133] = 8'hA2;
Memory[12132] = 8'h03;
Memory[12139] = 8'h00;
Memory[12138] = 8'h32;
Memory[12137] = 8'h22;
Memory[12136] = 8'hB3;
Memory[12143] = 8'h00;
Memory[12142] = 8'h02;
Memory[12141] = 8'h84;
Memory[12140] = 8'h63;
Memory[12147] = 8'h4E;
Memory[12146] = 8'h80;
Memory[12145] = 8'h50;
Memory[12144] = 8'h6F;
Memory[12151] = 8'h35;
Memory[12150] = 8'hCC;
Memory[12149] = 8'hA2;
Memory[12148] = 8'h03;
Memory[12155] = 8'h00;
Memory[12154] = 8'h32;
Memory[12153] = 8'h22;
Memory[12152] = 8'hB3;
Memory[12159] = 8'h00;
Memory[12158] = 8'h02;
Memory[12157] = 8'h84;
Memory[12156] = 8'h63;
Memory[12163] = 8'h4D;
Memory[12162] = 8'hC0;
Memory[12161] = 8'h50;
Memory[12160] = 8'h6F;
Memory[12167] = 8'h35;
Memory[12166] = 8'h8C;
Memory[12165] = 8'hA2;
Memory[12164] = 8'h03;
Memory[12171] = 8'h00;
Memory[12170] = 8'h32;
Memory[12169] = 8'h22;
Memory[12168] = 8'hB3;
Memory[12175] = 8'h00;
Memory[12174] = 8'h02;
Memory[12173] = 8'h84;
Memory[12172] = 8'h63;
Memory[12179] = 8'h4D;
Memory[12178] = 8'h00;
Memory[12177] = 8'h50;
Memory[12176] = 8'h6F;
Memory[12183] = 8'h35;
Memory[12182] = 8'h4C;
Memory[12181] = 8'hA2;
Memory[12180] = 8'h03;
Memory[12187] = 8'h00;
Memory[12186] = 8'h32;
Memory[12185] = 8'h22;
Memory[12184] = 8'hB3;
Memory[12191] = 8'h00;
Memory[12190] = 8'h02;
Memory[12189] = 8'h84;
Memory[12188] = 8'h63;
Memory[12195] = 8'h4C;
Memory[12194] = 8'h40;
Memory[12193] = 8'h50;
Memory[12192] = 8'h6F;
Memory[12199] = 8'h35;
Memory[12198] = 8'h0C;
Memory[12197] = 8'hA2;
Memory[12196] = 8'h03;
Memory[12203] = 8'h00;
Memory[12202] = 8'h32;
Memory[12201] = 8'h22;
Memory[12200] = 8'hB3;
Memory[12207] = 8'h00;
Memory[12206] = 8'h02;
Memory[12205] = 8'h84;
Memory[12204] = 8'h63;
Memory[12211] = 8'h4B;
Memory[12210] = 8'h80;
Memory[12209] = 8'h50;
Memory[12208] = 8'h6F;
Memory[12215] = 8'h34;
Memory[12214] = 8'hCC;
Memory[12213] = 8'hA2;
Memory[12212] = 8'h03;
Memory[12219] = 8'h00;
Memory[12218] = 8'h32;
Memory[12217] = 8'h22;
Memory[12216] = 8'hB3;
Memory[12223] = 8'h00;
Memory[12222] = 8'h02;
Memory[12221] = 8'h84;
Memory[12220] = 8'h63;
Memory[12227] = 8'h4A;
Memory[12226] = 8'hC0;
Memory[12225] = 8'h50;
Memory[12224] = 8'h6F;
Memory[12231] = 8'h34;
Memory[12230] = 8'h8C;
Memory[12229] = 8'hA2;
Memory[12228] = 8'h03;
Memory[12235] = 8'h00;
Memory[12234] = 8'h32;
Memory[12233] = 8'h22;
Memory[12232] = 8'hB3;
Memory[12239] = 8'h00;
Memory[12238] = 8'h02;
Memory[12237] = 8'h84;
Memory[12236] = 8'h63;
Memory[12243] = 8'h4A;
Memory[12242] = 8'h00;
Memory[12241] = 8'h50;
Memory[12240] = 8'h6F;
Memory[12247] = 8'h34;
Memory[12246] = 8'h4C;
Memory[12245] = 8'hA2;
Memory[12244] = 8'h03;
Memory[12251] = 8'h00;
Memory[12250] = 8'h32;
Memory[12249] = 8'h22;
Memory[12248] = 8'hB3;
Memory[12255] = 8'h00;
Memory[12254] = 8'h02;
Memory[12253] = 8'h84;
Memory[12252] = 8'h63;
Memory[12259] = 8'h49;
Memory[12258] = 8'h40;
Memory[12257] = 8'h50;
Memory[12256] = 8'h6F;
Memory[12263] = 8'h34;
Memory[12262] = 8'h0C;
Memory[12261] = 8'hA2;
Memory[12260] = 8'h03;
Memory[12267] = 8'h00;
Memory[12266] = 8'h32;
Memory[12265] = 8'h22;
Memory[12264] = 8'hB3;
Memory[12271] = 8'h00;
Memory[12270] = 8'h02;
Memory[12269] = 8'h84;
Memory[12268] = 8'h63;
Memory[12275] = 8'h48;
Memory[12274] = 8'h80;
Memory[12273] = 8'h50;
Memory[12272] = 8'h6F;
Memory[12279] = 8'h33;
Memory[12278] = 8'hCC;
Memory[12277] = 8'hA2;
Memory[12276] = 8'h03;
Memory[12283] = 8'h00;
Memory[12282] = 8'h32;
Memory[12281] = 8'h22;
Memory[12280] = 8'hB3;
Memory[12287] = 8'h00;
Memory[12286] = 8'h02;
Memory[12285] = 8'h84;
Memory[12284] = 8'h63;
Memory[12291] = 8'h47;
Memory[12290] = 8'hC0;
Memory[12289] = 8'h50;
Memory[12288] = 8'h6F;
Memory[12295] = 8'h33;
Memory[12294] = 8'h8C;
Memory[12293] = 8'hA2;
Memory[12292] = 8'h03;
Memory[12299] = 8'h00;
Memory[12298] = 8'h32;
Memory[12297] = 8'h22;
Memory[12296] = 8'hB3;
Memory[12303] = 8'h00;
Memory[12302] = 8'h02;
Memory[12301] = 8'h84;
Memory[12300] = 8'h63;
Memory[12307] = 8'h47;
Memory[12306] = 8'h00;
Memory[12305] = 8'h50;
Memory[12304] = 8'h6F;
Memory[12311] = 8'h33;
Memory[12310] = 8'h4C;
Memory[12309] = 8'hA2;
Memory[12308] = 8'h03;
Memory[12315] = 8'h00;
Memory[12314] = 8'h32;
Memory[12313] = 8'h22;
Memory[12312] = 8'hB3;
Memory[12319] = 8'h00;
Memory[12318] = 8'h02;
Memory[12317] = 8'h84;
Memory[12316] = 8'h63;
Memory[12323] = 8'h46;
Memory[12322] = 8'h40;
Memory[12321] = 8'h50;
Memory[12320] = 8'h6F;
Memory[12327] = 8'h33;
Memory[12326] = 8'h0C;
Memory[12325] = 8'hA2;
Memory[12324] = 8'h03;
Memory[12331] = 8'h00;
Memory[12330] = 8'h32;
Memory[12329] = 8'h22;
Memory[12328] = 8'hB3;
Memory[12335] = 8'h00;
Memory[12334] = 8'h02;
Memory[12333] = 8'h84;
Memory[12332] = 8'h63;
Memory[12339] = 8'h45;
Memory[12338] = 8'h80;
Memory[12337] = 8'h50;
Memory[12336] = 8'h6F;
Memory[12343] = 8'h32;
Memory[12342] = 8'hCC;
Memory[12341] = 8'hA2;
Memory[12340] = 8'h03;
Memory[12347] = 8'h00;
Memory[12346] = 8'h32;
Memory[12345] = 8'h22;
Memory[12344] = 8'hB3;
Memory[12351] = 8'h00;
Memory[12350] = 8'h02;
Memory[12349] = 8'h84;
Memory[12348] = 8'h63;
Memory[12355] = 8'h44;
Memory[12354] = 8'hC0;
Memory[12353] = 8'h50;
Memory[12352] = 8'h6F;
Memory[12359] = 8'h32;
Memory[12358] = 8'h8C;
Memory[12357] = 8'hA2;
Memory[12356] = 8'h03;
Memory[12363] = 8'h00;
Memory[12362] = 8'h32;
Memory[12361] = 8'h22;
Memory[12360] = 8'hB3;
Memory[12367] = 8'h00;
Memory[12366] = 8'h02;
Memory[12365] = 8'h84;
Memory[12364] = 8'h63;
Memory[12371] = 8'h44;
Memory[12370] = 8'h00;
Memory[12369] = 8'h50;
Memory[12368] = 8'h6F;
Memory[12375] = 8'h32;
Memory[12374] = 8'h4C;
Memory[12373] = 8'hA2;
Memory[12372] = 8'h03;
Memory[12379] = 8'h00;
Memory[12378] = 8'h32;
Memory[12377] = 8'h22;
Memory[12376] = 8'hB3;
Memory[12383] = 8'h00;
Memory[12382] = 8'h02;
Memory[12381] = 8'h84;
Memory[12380] = 8'h63;
Memory[12387] = 8'h43;
Memory[12386] = 8'h40;
Memory[12385] = 8'h50;
Memory[12384] = 8'h6F;
Memory[12391] = 8'h32;
Memory[12390] = 8'h0C;
Memory[12389] = 8'hA2;
Memory[12388] = 8'h03;
Memory[12395] = 8'h00;
Memory[12394] = 8'h32;
Memory[12393] = 8'h22;
Memory[12392] = 8'hB3;
Memory[12399] = 8'h00;
Memory[12398] = 8'h02;
Memory[12397] = 8'h84;
Memory[12396] = 8'h63;
Memory[12403] = 8'h42;
Memory[12402] = 8'h80;
Memory[12401] = 8'h50;
Memory[12400] = 8'h6F;
Memory[12407] = 8'h31;
Memory[12406] = 8'hCC;
Memory[12405] = 8'hA2;
Memory[12404] = 8'h03;
Memory[12411] = 8'h00;
Memory[12410] = 8'h32;
Memory[12409] = 8'h22;
Memory[12408] = 8'hB3;
Memory[12415] = 8'h00;
Memory[12414] = 8'h02;
Memory[12413] = 8'h84;
Memory[12412] = 8'h63;
Memory[12419] = 8'h41;
Memory[12418] = 8'hC0;
Memory[12417] = 8'h50;
Memory[12416] = 8'h6F;
Memory[12423] = 8'h31;
Memory[12422] = 8'h8C;
Memory[12421] = 8'hA2;
Memory[12420] = 8'h03;
Memory[12427] = 8'h00;
Memory[12426] = 8'h32;
Memory[12425] = 8'h22;
Memory[12424] = 8'hB3;
Memory[12431] = 8'h00;
Memory[12430] = 8'h02;
Memory[12429] = 8'h84;
Memory[12428] = 8'h63;
Memory[12435] = 8'h41;
Memory[12434] = 8'h00;
Memory[12433] = 8'h50;
Memory[12432] = 8'h6F;
Memory[12439] = 8'h31;
Memory[12438] = 8'h4C;
Memory[12437] = 8'hA2;
Memory[12436] = 8'h03;
Memory[12443] = 8'h00;
Memory[12442] = 8'h32;
Memory[12441] = 8'h22;
Memory[12440] = 8'hB3;
Memory[12447] = 8'h00;
Memory[12446] = 8'h02;
Memory[12445] = 8'h84;
Memory[12444] = 8'h63;
Memory[12451] = 8'h40;
Memory[12450] = 8'h40;
Memory[12449] = 8'h50;
Memory[12448] = 8'h6F;
Memory[12455] = 8'h31;
Memory[12454] = 8'h0C;
Memory[12453] = 8'hA2;
Memory[12452] = 8'h03;
Memory[12459] = 8'h00;
Memory[12458] = 8'h32;
Memory[12457] = 8'h22;
Memory[12456] = 8'hB3;
Memory[12463] = 8'h00;
Memory[12462] = 8'h02;
Memory[12461] = 8'h84;
Memory[12460] = 8'h63;
Memory[12467] = 8'h3F;
Memory[12466] = 8'h80;
Memory[12465] = 8'h50;
Memory[12464] = 8'h6F;
Memory[12471] = 8'h30;
Memory[12470] = 8'hCC;
Memory[12469] = 8'hA2;
Memory[12468] = 8'h03;
Memory[12475] = 8'h00;
Memory[12474] = 8'h32;
Memory[12473] = 8'h22;
Memory[12472] = 8'hB3;
Memory[12479] = 8'h00;
Memory[12478] = 8'h02;
Memory[12477] = 8'h84;
Memory[12476] = 8'h63;
Memory[12483] = 8'h3E;
Memory[12482] = 8'hC0;
Memory[12481] = 8'h50;
Memory[12480] = 8'h6F;
Memory[12487] = 8'h30;
Memory[12486] = 8'h8C;
Memory[12485] = 8'hA2;
Memory[12484] = 8'h03;
Memory[12491] = 8'h00;
Memory[12490] = 8'h32;
Memory[12489] = 8'h22;
Memory[12488] = 8'hB3;
Memory[12495] = 8'h00;
Memory[12494] = 8'h02;
Memory[12493] = 8'h84;
Memory[12492] = 8'h63;
Memory[12499] = 8'h3E;
Memory[12498] = 8'h00;
Memory[12497] = 8'h50;
Memory[12496] = 8'h6F;
Memory[12503] = 8'h30;
Memory[12502] = 8'h4C;
Memory[12501] = 8'hA2;
Memory[12500] = 8'h03;
Memory[12507] = 8'h00;
Memory[12506] = 8'h32;
Memory[12505] = 8'h22;
Memory[12504] = 8'hB3;
Memory[12511] = 8'h00;
Memory[12510] = 8'h02;
Memory[12509] = 8'h84;
Memory[12508] = 8'h63;
Memory[12515] = 8'h3D;
Memory[12514] = 8'h40;
Memory[12513] = 8'h50;
Memory[12512] = 8'h6F;
Memory[12519] = 8'h30;
Memory[12518] = 8'h0C;
Memory[12517] = 8'hA2;
Memory[12516] = 8'h03;
Memory[12523] = 8'h00;
Memory[12522] = 8'h32;
Memory[12521] = 8'h22;
Memory[12520] = 8'hB3;
Memory[12527] = 8'h00;
Memory[12526] = 8'h02;
Memory[12525] = 8'h84;
Memory[12524] = 8'h63;
Memory[12531] = 8'h3C;
Memory[12530] = 8'h80;
Memory[12529] = 8'h50;
Memory[12528] = 8'h6F;
Memory[12535] = 8'h2F;
Memory[12534] = 8'hCC;
Memory[12533] = 8'hA2;
Memory[12532] = 8'h03;
Memory[12539] = 8'h00;
Memory[12538] = 8'h32;
Memory[12537] = 8'h22;
Memory[12536] = 8'hB3;
Memory[12543] = 8'h00;
Memory[12542] = 8'h02;
Memory[12541] = 8'h84;
Memory[12540] = 8'h63;
Memory[12547] = 8'h3B;
Memory[12546] = 8'hC0;
Memory[12545] = 8'h50;
Memory[12544] = 8'h6F;
Memory[12551] = 8'h2F;
Memory[12550] = 8'h8C;
Memory[12549] = 8'hA2;
Memory[12548] = 8'h03;
Memory[12555] = 8'h00;
Memory[12554] = 8'h32;
Memory[12553] = 8'h22;
Memory[12552] = 8'hB3;
Memory[12559] = 8'h00;
Memory[12558] = 8'h02;
Memory[12557] = 8'h84;
Memory[12556] = 8'h63;
Memory[12563] = 8'h3B;
Memory[12562] = 8'h00;
Memory[12561] = 8'h50;
Memory[12560] = 8'h6F;
Memory[12567] = 8'h2F;
Memory[12566] = 8'h4C;
Memory[12565] = 8'hA2;
Memory[12564] = 8'h03;
Memory[12571] = 8'h00;
Memory[12570] = 8'h32;
Memory[12569] = 8'h22;
Memory[12568] = 8'hB3;
Memory[12575] = 8'h00;
Memory[12574] = 8'h02;
Memory[12573] = 8'h84;
Memory[12572] = 8'h63;
Memory[12579] = 8'h3A;
Memory[12578] = 8'h40;
Memory[12577] = 8'h50;
Memory[12576] = 8'h6F;
Memory[12583] = 8'h2F;
Memory[12582] = 8'h0C;
Memory[12581] = 8'hA2;
Memory[12580] = 8'h03;
Memory[12587] = 8'h00;
Memory[12586] = 8'h32;
Memory[12585] = 8'h22;
Memory[12584] = 8'hB3;
Memory[12591] = 8'h00;
Memory[12590] = 8'h02;
Memory[12589] = 8'h84;
Memory[12588] = 8'h63;
Memory[12595] = 8'h39;
Memory[12594] = 8'h80;
Memory[12593] = 8'h50;
Memory[12592] = 8'h6F;
Memory[12599] = 8'h2E;
Memory[12598] = 8'hCC;
Memory[12597] = 8'hA2;
Memory[12596] = 8'h03;
Memory[12603] = 8'h00;
Memory[12602] = 8'h32;
Memory[12601] = 8'h22;
Memory[12600] = 8'hB3;
Memory[12607] = 8'h00;
Memory[12606] = 8'h02;
Memory[12605] = 8'h84;
Memory[12604] = 8'h63;
Memory[12611] = 8'h38;
Memory[12610] = 8'hC0;
Memory[12609] = 8'h50;
Memory[12608] = 8'h6F;
Memory[12615] = 8'h2E;
Memory[12614] = 8'h8C;
Memory[12613] = 8'hA2;
Memory[12612] = 8'h03;
Memory[12619] = 8'h00;
Memory[12618] = 8'h32;
Memory[12617] = 8'h22;
Memory[12616] = 8'hB3;
Memory[12623] = 8'h00;
Memory[12622] = 8'h02;
Memory[12621] = 8'h84;
Memory[12620] = 8'h63;
Memory[12627] = 8'h38;
Memory[12626] = 8'h00;
Memory[12625] = 8'h50;
Memory[12624] = 8'h6F;
Memory[12631] = 8'h2E;
Memory[12630] = 8'h4C;
Memory[12629] = 8'hA2;
Memory[12628] = 8'h03;
Memory[12635] = 8'h00;
Memory[12634] = 8'h32;
Memory[12633] = 8'h22;
Memory[12632] = 8'hB3;
Memory[12639] = 8'h00;
Memory[12638] = 8'h02;
Memory[12637] = 8'h84;
Memory[12636] = 8'h63;
Memory[12643] = 8'h37;
Memory[12642] = 8'h40;
Memory[12641] = 8'h50;
Memory[12640] = 8'h6F;
Memory[12647] = 8'h2E;
Memory[12646] = 8'h0C;
Memory[12645] = 8'hA2;
Memory[12644] = 8'h03;
Memory[12651] = 8'h00;
Memory[12650] = 8'h32;
Memory[12649] = 8'h22;
Memory[12648] = 8'hB3;
Memory[12655] = 8'h00;
Memory[12654] = 8'h02;
Memory[12653] = 8'h84;
Memory[12652] = 8'h63;
Memory[12659] = 8'h36;
Memory[12658] = 8'h80;
Memory[12657] = 8'h50;
Memory[12656] = 8'h6F;
Memory[12663] = 8'h2D;
Memory[12662] = 8'hCC;
Memory[12661] = 8'hA2;
Memory[12660] = 8'h03;
Memory[12667] = 8'h00;
Memory[12666] = 8'h32;
Memory[12665] = 8'h22;
Memory[12664] = 8'hB3;
Memory[12671] = 8'h00;
Memory[12670] = 8'h02;
Memory[12669] = 8'h84;
Memory[12668] = 8'h63;
Memory[12675] = 8'h35;
Memory[12674] = 8'hC0;
Memory[12673] = 8'h50;
Memory[12672] = 8'h6F;
Memory[12679] = 8'h2D;
Memory[12678] = 8'h8C;
Memory[12677] = 8'hA2;
Memory[12676] = 8'h03;
Memory[12683] = 8'h00;
Memory[12682] = 8'h32;
Memory[12681] = 8'h22;
Memory[12680] = 8'hB3;
Memory[12687] = 8'h00;
Memory[12686] = 8'h02;
Memory[12685] = 8'h84;
Memory[12684] = 8'h63;
Memory[12691] = 8'h35;
Memory[12690] = 8'h00;
Memory[12689] = 8'h50;
Memory[12688] = 8'h6F;
Memory[12695] = 8'h2D;
Memory[12694] = 8'h4C;
Memory[12693] = 8'hA2;
Memory[12692] = 8'h03;
Memory[12699] = 8'h00;
Memory[12698] = 8'h32;
Memory[12697] = 8'h22;
Memory[12696] = 8'hB3;
Memory[12703] = 8'h00;
Memory[12702] = 8'h02;
Memory[12701] = 8'h84;
Memory[12700] = 8'h63;
Memory[12707] = 8'h34;
Memory[12706] = 8'h40;
Memory[12705] = 8'h50;
Memory[12704] = 8'h6F;
Memory[12711] = 8'h2D;
Memory[12710] = 8'h0C;
Memory[12709] = 8'hA2;
Memory[12708] = 8'h03;
Memory[12715] = 8'h00;
Memory[12714] = 8'h32;
Memory[12713] = 8'h22;
Memory[12712] = 8'hB3;
Memory[12719] = 8'h00;
Memory[12718] = 8'h02;
Memory[12717] = 8'h84;
Memory[12716] = 8'h63;
Memory[12723] = 8'h33;
Memory[12722] = 8'h80;
Memory[12721] = 8'h50;
Memory[12720] = 8'h6F;
Memory[12727] = 8'h2C;
Memory[12726] = 8'hCC;
Memory[12725] = 8'hA2;
Memory[12724] = 8'h03;
Memory[12731] = 8'h00;
Memory[12730] = 8'h32;
Memory[12729] = 8'h22;
Memory[12728] = 8'hB3;
Memory[12735] = 8'h00;
Memory[12734] = 8'h02;
Memory[12733] = 8'h84;
Memory[12732] = 8'h63;
Memory[12739] = 8'h32;
Memory[12738] = 8'hC0;
Memory[12737] = 8'h50;
Memory[12736] = 8'h6F;
Memory[12743] = 8'h2C;
Memory[12742] = 8'h8C;
Memory[12741] = 8'hA2;
Memory[12740] = 8'h03;
Memory[12747] = 8'h00;
Memory[12746] = 8'h32;
Memory[12745] = 8'h22;
Memory[12744] = 8'hB3;
Memory[12751] = 8'h00;
Memory[12750] = 8'h02;
Memory[12749] = 8'h84;
Memory[12748] = 8'h63;
Memory[12755] = 8'h32;
Memory[12754] = 8'h00;
Memory[12753] = 8'h50;
Memory[12752] = 8'h6F;
Memory[12759] = 8'h2C;
Memory[12758] = 8'h4C;
Memory[12757] = 8'hA2;
Memory[12756] = 8'h03;
Memory[12763] = 8'h00;
Memory[12762] = 8'h32;
Memory[12761] = 8'h22;
Memory[12760] = 8'hB3;
Memory[12767] = 8'h00;
Memory[12766] = 8'h02;
Memory[12765] = 8'h84;
Memory[12764] = 8'h63;
Memory[12771] = 8'h31;
Memory[12770] = 8'h40;
Memory[12769] = 8'h50;
Memory[12768] = 8'h6F;
Memory[12775] = 8'h2C;
Memory[12774] = 8'h0C;
Memory[12773] = 8'hA2;
Memory[12772] = 8'h03;
Memory[12779] = 8'h00;
Memory[12778] = 8'h32;
Memory[12777] = 8'h22;
Memory[12776] = 8'hB3;
Memory[12783] = 8'h00;
Memory[12782] = 8'h02;
Memory[12781] = 8'h84;
Memory[12780] = 8'h63;
Memory[12787] = 8'h30;
Memory[12786] = 8'h80;
Memory[12785] = 8'h50;
Memory[12784] = 8'h6F;
Memory[12791] = 8'h2B;
Memory[12790] = 8'hCC;
Memory[12789] = 8'hA2;
Memory[12788] = 8'h03;
Memory[12795] = 8'h00;
Memory[12794] = 8'h32;
Memory[12793] = 8'h22;
Memory[12792] = 8'hB3;
Memory[12799] = 8'h00;
Memory[12798] = 8'h02;
Memory[12797] = 8'h84;
Memory[12796] = 8'h63;
Memory[12803] = 8'h2F;
Memory[12802] = 8'hC0;
Memory[12801] = 8'h50;
Memory[12800] = 8'h6F;
Memory[12807] = 8'h2B;
Memory[12806] = 8'h8C;
Memory[12805] = 8'hA2;
Memory[12804] = 8'h03;
Memory[12811] = 8'h00;
Memory[12810] = 8'h32;
Memory[12809] = 8'h22;
Memory[12808] = 8'hB3;
Memory[12815] = 8'h00;
Memory[12814] = 8'h02;
Memory[12813] = 8'h84;
Memory[12812] = 8'h63;
Memory[12819] = 8'h2F;
Memory[12818] = 8'h00;
Memory[12817] = 8'h50;
Memory[12816] = 8'h6F;
Memory[12823] = 8'h2B;
Memory[12822] = 8'h4C;
Memory[12821] = 8'hA2;
Memory[12820] = 8'h03;
Memory[12827] = 8'h00;
Memory[12826] = 8'h32;
Memory[12825] = 8'h22;
Memory[12824] = 8'hB3;
Memory[12831] = 8'h00;
Memory[12830] = 8'h02;
Memory[12829] = 8'h84;
Memory[12828] = 8'h63;
Memory[12835] = 8'h2E;
Memory[12834] = 8'h40;
Memory[12833] = 8'h50;
Memory[12832] = 8'h6F;
Memory[12839] = 8'h2B;
Memory[12838] = 8'h0C;
Memory[12837] = 8'hA2;
Memory[12836] = 8'h03;
Memory[12843] = 8'h00;
Memory[12842] = 8'h32;
Memory[12841] = 8'h22;
Memory[12840] = 8'hB3;
Memory[12847] = 8'h00;
Memory[12846] = 8'h02;
Memory[12845] = 8'h84;
Memory[12844] = 8'h63;
Memory[12851] = 8'h2D;
Memory[12850] = 8'h80;
Memory[12849] = 8'h50;
Memory[12848] = 8'h6F;
Memory[12855] = 8'h2A;
Memory[12854] = 8'hCC;
Memory[12853] = 8'hA2;
Memory[12852] = 8'h03;
Memory[12859] = 8'h00;
Memory[12858] = 8'h32;
Memory[12857] = 8'h22;
Memory[12856] = 8'hB3;
Memory[12863] = 8'h00;
Memory[12862] = 8'h02;
Memory[12861] = 8'h84;
Memory[12860] = 8'h63;
Memory[12867] = 8'h2C;
Memory[12866] = 8'hC0;
Memory[12865] = 8'h50;
Memory[12864] = 8'h6F;
Memory[12871] = 8'h2A;
Memory[12870] = 8'h8C;
Memory[12869] = 8'hA2;
Memory[12868] = 8'h03;
Memory[12875] = 8'h00;
Memory[12874] = 8'h32;
Memory[12873] = 8'h22;
Memory[12872] = 8'hB3;
Memory[12879] = 8'h00;
Memory[12878] = 8'h02;
Memory[12877] = 8'h84;
Memory[12876] = 8'h63;
Memory[12883] = 8'h2C;
Memory[12882] = 8'h00;
Memory[12881] = 8'h50;
Memory[12880] = 8'h6F;
Memory[12887] = 8'h2A;
Memory[12886] = 8'h4C;
Memory[12885] = 8'hA2;
Memory[12884] = 8'h03;
Memory[12891] = 8'h00;
Memory[12890] = 8'h32;
Memory[12889] = 8'h22;
Memory[12888] = 8'hB3;
Memory[12895] = 8'h00;
Memory[12894] = 8'h02;
Memory[12893] = 8'h84;
Memory[12892] = 8'h63;
Memory[12899] = 8'h2B;
Memory[12898] = 8'h40;
Memory[12897] = 8'h50;
Memory[12896] = 8'h6F;
Memory[12903] = 8'h2A;
Memory[12902] = 8'h0C;
Memory[12901] = 8'hA2;
Memory[12900] = 8'h03;
Memory[12907] = 8'h00;
Memory[12906] = 8'h32;
Memory[12905] = 8'h22;
Memory[12904] = 8'hB3;
Memory[12911] = 8'h00;
Memory[12910] = 8'h02;
Memory[12909] = 8'h84;
Memory[12908] = 8'h63;
Memory[12915] = 8'h2A;
Memory[12914] = 8'h80;
Memory[12913] = 8'h50;
Memory[12912] = 8'h6F;
Memory[12919] = 8'h29;
Memory[12918] = 8'hCC;
Memory[12917] = 8'hA2;
Memory[12916] = 8'h03;
Memory[12923] = 8'h00;
Memory[12922] = 8'h32;
Memory[12921] = 8'h22;
Memory[12920] = 8'hB3;
Memory[12927] = 8'h00;
Memory[12926] = 8'h02;
Memory[12925] = 8'h84;
Memory[12924] = 8'h63;
Memory[12931] = 8'h29;
Memory[12930] = 8'hC0;
Memory[12929] = 8'h50;
Memory[12928] = 8'h6F;
Memory[12935] = 8'h29;
Memory[12934] = 8'h8C;
Memory[12933] = 8'hA2;
Memory[12932] = 8'h03;
Memory[12939] = 8'h00;
Memory[12938] = 8'h32;
Memory[12937] = 8'h22;
Memory[12936] = 8'hB3;
Memory[12943] = 8'h00;
Memory[12942] = 8'h02;
Memory[12941] = 8'h84;
Memory[12940] = 8'h63;
Memory[12947] = 8'h29;
Memory[12946] = 8'h00;
Memory[12945] = 8'h50;
Memory[12944] = 8'h6F;
Memory[12951] = 8'h29;
Memory[12950] = 8'h4C;
Memory[12949] = 8'hA2;
Memory[12948] = 8'h03;
Memory[12955] = 8'h00;
Memory[12954] = 8'h32;
Memory[12953] = 8'h22;
Memory[12952] = 8'hB3;
Memory[12959] = 8'h00;
Memory[12958] = 8'h02;
Memory[12957] = 8'h84;
Memory[12956] = 8'h63;
Memory[12963] = 8'h28;
Memory[12962] = 8'h40;
Memory[12961] = 8'h50;
Memory[12960] = 8'h6F;
Memory[12967] = 8'h29;
Memory[12966] = 8'h0C;
Memory[12965] = 8'hA2;
Memory[12964] = 8'h03;
Memory[12971] = 8'h00;
Memory[12970] = 8'h32;
Memory[12969] = 8'h22;
Memory[12968] = 8'hB3;
Memory[12975] = 8'h00;
Memory[12974] = 8'h02;
Memory[12973] = 8'h84;
Memory[12972] = 8'h63;
Memory[12979] = 8'h27;
Memory[12978] = 8'h80;
Memory[12977] = 8'h50;
Memory[12976] = 8'h6F;
Memory[12983] = 8'h28;
Memory[12982] = 8'hCC;
Memory[12981] = 8'hA2;
Memory[12980] = 8'h03;
Memory[12987] = 8'h00;
Memory[12986] = 8'h32;
Memory[12985] = 8'h22;
Memory[12984] = 8'hB3;
Memory[12991] = 8'h00;
Memory[12990] = 8'h02;
Memory[12989] = 8'h84;
Memory[12988] = 8'h63;
Memory[12995] = 8'h26;
Memory[12994] = 8'hC0;
Memory[12993] = 8'h50;
Memory[12992] = 8'h6F;
Memory[12999] = 8'h28;
Memory[12998] = 8'h8C;
Memory[12997] = 8'hA2;
Memory[12996] = 8'h03;
Memory[13003] = 8'h00;
Memory[13002] = 8'h32;
Memory[13001] = 8'h22;
Memory[13000] = 8'hB3;
Memory[13007] = 8'h00;
Memory[13006] = 8'h02;
Memory[13005] = 8'h84;
Memory[13004] = 8'h63;
Memory[13011] = 8'h26;
Memory[13010] = 8'h00;
Memory[13009] = 8'h50;
Memory[13008] = 8'h6F;
Memory[13015] = 8'h28;
Memory[13014] = 8'h4C;
Memory[13013] = 8'hA2;
Memory[13012] = 8'h03;
Memory[13019] = 8'h00;
Memory[13018] = 8'h32;
Memory[13017] = 8'h22;
Memory[13016] = 8'hB3;
Memory[13023] = 8'h00;
Memory[13022] = 8'h02;
Memory[13021] = 8'h84;
Memory[13020] = 8'h63;
Memory[13027] = 8'h25;
Memory[13026] = 8'h40;
Memory[13025] = 8'h50;
Memory[13024] = 8'h6F;
Memory[13031] = 8'h28;
Memory[13030] = 8'h0C;
Memory[13029] = 8'hA2;
Memory[13028] = 8'h03;
Memory[13035] = 8'h00;
Memory[13034] = 8'h32;
Memory[13033] = 8'h22;
Memory[13032] = 8'hB3;
Memory[13039] = 8'h00;
Memory[13038] = 8'h02;
Memory[13037] = 8'h84;
Memory[13036] = 8'h63;
Memory[13043] = 8'h24;
Memory[13042] = 8'h80;
Memory[13041] = 8'h50;
Memory[13040] = 8'h6F;
Memory[13047] = 8'h27;
Memory[13046] = 8'hCC;
Memory[13045] = 8'hA2;
Memory[13044] = 8'h03;
Memory[13051] = 8'h00;
Memory[13050] = 8'h32;
Memory[13049] = 8'h22;
Memory[13048] = 8'hB3;
Memory[13055] = 8'h00;
Memory[13054] = 8'h02;
Memory[13053] = 8'h84;
Memory[13052] = 8'h63;
Memory[13059] = 8'h23;
Memory[13058] = 8'hC0;
Memory[13057] = 8'h50;
Memory[13056] = 8'h6F;
Memory[13063] = 8'h27;
Memory[13062] = 8'h8C;
Memory[13061] = 8'hA2;
Memory[13060] = 8'h03;
Memory[13067] = 8'h00;
Memory[13066] = 8'h32;
Memory[13065] = 8'h22;
Memory[13064] = 8'hB3;
Memory[13071] = 8'h00;
Memory[13070] = 8'h02;
Memory[13069] = 8'h84;
Memory[13068] = 8'h63;
Memory[13075] = 8'h23;
Memory[13074] = 8'h00;
Memory[13073] = 8'h50;
Memory[13072] = 8'h6F;
Memory[13079] = 8'h27;
Memory[13078] = 8'h4C;
Memory[13077] = 8'hA2;
Memory[13076] = 8'h03;
Memory[13083] = 8'h00;
Memory[13082] = 8'h32;
Memory[13081] = 8'h22;
Memory[13080] = 8'hB3;
Memory[13087] = 8'h00;
Memory[13086] = 8'h02;
Memory[13085] = 8'h84;
Memory[13084] = 8'h63;
Memory[13091] = 8'h22;
Memory[13090] = 8'h40;
Memory[13089] = 8'h50;
Memory[13088] = 8'h6F;
Memory[13095] = 8'h27;
Memory[13094] = 8'h0C;
Memory[13093] = 8'hA2;
Memory[13092] = 8'h03;
Memory[13099] = 8'h00;
Memory[13098] = 8'h32;
Memory[13097] = 8'h22;
Memory[13096] = 8'hB3;
Memory[13103] = 8'h00;
Memory[13102] = 8'h02;
Memory[13101] = 8'h84;
Memory[13100] = 8'h63;
Memory[13107] = 8'h21;
Memory[13106] = 8'h80;
Memory[13105] = 8'h50;
Memory[13104] = 8'h6F;
Memory[13111] = 8'h26;
Memory[13110] = 8'hCC;
Memory[13109] = 8'hA2;
Memory[13108] = 8'h03;
Memory[13115] = 8'h00;
Memory[13114] = 8'h32;
Memory[13113] = 8'h22;
Memory[13112] = 8'hB3;
Memory[13119] = 8'h00;
Memory[13118] = 8'h02;
Memory[13117] = 8'h84;
Memory[13116] = 8'h63;
Memory[13123] = 8'h20;
Memory[13122] = 8'hC0;
Memory[13121] = 8'h50;
Memory[13120] = 8'h6F;
Memory[13127] = 8'h26;
Memory[13126] = 8'h8C;
Memory[13125] = 8'hA2;
Memory[13124] = 8'h03;
Memory[13131] = 8'h00;
Memory[13130] = 8'h32;
Memory[13129] = 8'h22;
Memory[13128] = 8'hB3;
Memory[13135] = 8'h00;
Memory[13134] = 8'h02;
Memory[13133] = 8'h84;
Memory[13132] = 8'h63;
Memory[13139] = 8'h20;
Memory[13138] = 8'h00;
Memory[13137] = 8'h50;
Memory[13136] = 8'h6F;
Memory[13143] = 8'h26;
Memory[13142] = 8'h4C;
Memory[13141] = 8'hA2;
Memory[13140] = 8'h03;
Memory[13147] = 8'h00;
Memory[13146] = 8'h32;
Memory[13145] = 8'h22;
Memory[13144] = 8'hB3;
Memory[13151] = 8'h00;
Memory[13150] = 8'h02;
Memory[13149] = 8'h84;
Memory[13148] = 8'h63;
Memory[13155] = 8'h1F;
Memory[13154] = 8'h40;
Memory[13153] = 8'h50;
Memory[13152] = 8'h6F;
Memory[13159] = 8'h26;
Memory[13158] = 8'h0C;
Memory[13157] = 8'hA2;
Memory[13156] = 8'h03;
Memory[13163] = 8'h00;
Memory[13162] = 8'h32;
Memory[13161] = 8'h22;
Memory[13160] = 8'hB3;
Memory[13167] = 8'h00;
Memory[13166] = 8'h02;
Memory[13165] = 8'h84;
Memory[13164] = 8'h63;
Memory[13171] = 8'h1E;
Memory[13170] = 8'h80;
Memory[13169] = 8'h50;
Memory[13168] = 8'h6F;
Memory[13175] = 8'h25;
Memory[13174] = 8'hCC;
Memory[13173] = 8'hA2;
Memory[13172] = 8'h03;
Memory[13179] = 8'h00;
Memory[13178] = 8'h32;
Memory[13177] = 8'h22;
Memory[13176] = 8'hB3;
Memory[13183] = 8'h00;
Memory[13182] = 8'h02;
Memory[13181] = 8'h84;
Memory[13180] = 8'h63;
Memory[13187] = 8'h1D;
Memory[13186] = 8'hC0;
Memory[13185] = 8'h50;
Memory[13184] = 8'h6F;
Memory[13191] = 8'h25;
Memory[13190] = 8'h8C;
Memory[13189] = 8'hA2;
Memory[13188] = 8'h03;
Memory[13195] = 8'h00;
Memory[13194] = 8'h32;
Memory[13193] = 8'h22;
Memory[13192] = 8'hB3;
Memory[13199] = 8'h00;
Memory[13198] = 8'h02;
Memory[13197] = 8'h84;
Memory[13196] = 8'h63;
Memory[13203] = 8'h1D;
Memory[13202] = 8'h00;
Memory[13201] = 8'h50;
Memory[13200] = 8'h6F;
Memory[13207] = 8'h25;
Memory[13206] = 8'h4C;
Memory[13205] = 8'hA2;
Memory[13204] = 8'h03;
Memory[13211] = 8'h00;
Memory[13210] = 8'h32;
Memory[13209] = 8'h22;
Memory[13208] = 8'hB3;
Memory[13215] = 8'h00;
Memory[13214] = 8'h02;
Memory[13213] = 8'h84;
Memory[13212] = 8'h63;
Memory[13219] = 8'h1C;
Memory[13218] = 8'h40;
Memory[13217] = 8'h50;
Memory[13216] = 8'h6F;
Memory[13223] = 8'h25;
Memory[13222] = 8'h0C;
Memory[13221] = 8'hA2;
Memory[13220] = 8'h03;
Memory[13227] = 8'h00;
Memory[13226] = 8'h32;
Memory[13225] = 8'h22;
Memory[13224] = 8'hB3;
Memory[13231] = 8'h00;
Memory[13230] = 8'h02;
Memory[13229] = 8'h84;
Memory[13228] = 8'h63;
Memory[13235] = 8'h1B;
Memory[13234] = 8'h80;
Memory[13233] = 8'h50;
Memory[13232] = 8'h6F;
Memory[13239] = 8'h24;
Memory[13238] = 8'hCC;
Memory[13237] = 8'hA2;
Memory[13236] = 8'h03;
Memory[13243] = 8'h00;
Memory[13242] = 8'h32;
Memory[13241] = 8'h22;
Memory[13240] = 8'hB3;
Memory[13247] = 8'h00;
Memory[13246] = 8'h02;
Memory[13245] = 8'h84;
Memory[13244] = 8'h63;
Memory[13251] = 8'h1A;
Memory[13250] = 8'hC0;
Memory[13249] = 8'h50;
Memory[13248] = 8'h6F;
Memory[13255] = 8'h24;
Memory[13254] = 8'h8C;
Memory[13253] = 8'hA2;
Memory[13252] = 8'h03;
Memory[13259] = 8'h00;
Memory[13258] = 8'h32;
Memory[13257] = 8'h22;
Memory[13256] = 8'hB3;
Memory[13263] = 8'h00;
Memory[13262] = 8'h02;
Memory[13261] = 8'h84;
Memory[13260] = 8'h63;
Memory[13267] = 8'h1A;
Memory[13266] = 8'h00;
Memory[13265] = 8'h50;
Memory[13264] = 8'h6F;
Memory[13271] = 8'h24;
Memory[13270] = 8'h4C;
Memory[13269] = 8'hA2;
Memory[13268] = 8'h03;
Memory[13275] = 8'h00;
Memory[13274] = 8'h32;
Memory[13273] = 8'h22;
Memory[13272] = 8'hB3;
Memory[13279] = 8'h00;
Memory[13278] = 8'h02;
Memory[13277] = 8'h84;
Memory[13276] = 8'h63;
Memory[13283] = 8'h19;
Memory[13282] = 8'h40;
Memory[13281] = 8'h50;
Memory[13280] = 8'h6F;
Memory[13287] = 8'h24;
Memory[13286] = 8'h0C;
Memory[13285] = 8'hA2;
Memory[13284] = 8'h03;
Memory[13291] = 8'h00;
Memory[13290] = 8'h32;
Memory[13289] = 8'h22;
Memory[13288] = 8'hB3;
Memory[13295] = 8'h00;
Memory[13294] = 8'h02;
Memory[13293] = 8'h84;
Memory[13292] = 8'h63;
Memory[13299] = 8'h18;
Memory[13298] = 8'h80;
Memory[13297] = 8'h50;
Memory[13296] = 8'h6F;
Memory[13303] = 8'h23;
Memory[13302] = 8'hCC;
Memory[13301] = 8'hA2;
Memory[13300] = 8'h03;
Memory[13307] = 8'h00;
Memory[13306] = 8'h32;
Memory[13305] = 8'h22;
Memory[13304] = 8'hB3;
Memory[13311] = 8'h00;
Memory[13310] = 8'h02;
Memory[13309] = 8'h84;
Memory[13308] = 8'h63;
Memory[13315] = 8'h17;
Memory[13314] = 8'hC0;
Memory[13313] = 8'h50;
Memory[13312] = 8'h6F;
Memory[13319] = 8'h23;
Memory[13318] = 8'h8C;
Memory[13317] = 8'hA2;
Memory[13316] = 8'h03;
Memory[13323] = 8'h00;
Memory[13322] = 8'h32;
Memory[13321] = 8'h22;
Memory[13320] = 8'hB3;
Memory[13327] = 8'h00;
Memory[13326] = 8'h02;
Memory[13325] = 8'h84;
Memory[13324] = 8'h63;
Memory[13331] = 8'h17;
Memory[13330] = 8'h00;
Memory[13329] = 8'h50;
Memory[13328] = 8'h6F;
Memory[13335] = 8'h23;
Memory[13334] = 8'h4C;
Memory[13333] = 8'hA2;
Memory[13332] = 8'h03;
Memory[13339] = 8'h00;
Memory[13338] = 8'h32;
Memory[13337] = 8'h22;
Memory[13336] = 8'hB3;
Memory[13343] = 8'h00;
Memory[13342] = 8'h02;
Memory[13341] = 8'h84;
Memory[13340] = 8'h63;
Memory[13347] = 8'h16;
Memory[13346] = 8'h40;
Memory[13345] = 8'h50;
Memory[13344] = 8'h6F;
Memory[13351] = 8'h23;
Memory[13350] = 8'h0C;
Memory[13349] = 8'hA2;
Memory[13348] = 8'h03;
Memory[13355] = 8'h00;
Memory[13354] = 8'h32;
Memory[13353] = 8'h22;
Memory[13352] = 8'hB3;
Memory[13359] = 8'h00;
Memory[13358] = 8'h02;
Memory[13357] = 8'h84;
Memory[13356] = 8'h63;
Memory[13363] = 8'h15;
Memory[13362] = 8'h80;
Memory[13361] = 8'h50;
Memory[13360] = 8'h6F;
Memory[13367] = 8'h22;
Memory[13366] = 8'hCC;
Memory[13365] = 8'hA2;
Memory[13364] = 8'h03;
Memory[13371] = 8'h00;
Memory[13370] = 8'h32;
Memory[13369] = 8'h22;
Memory[13368] = 8'hB3;
Memory[13375] = 8'h00;
Memory[13374] = 8'h02;
Memory[13373] = 8'h84;
Memory[13372] = 8'h63;
Memory[13379] = 8'h14;
Memory[13378] = 8'hC0;
Memory[13377] = 8'h50;
Memory[13376] = 8'h6F;
Memory[13383] = 8'h22;
Memory[13382] = 8'h8C;
Memory[13381] = 8'hA2;
Memory[13380] = 8'h03;
Memory[13387] = 8'h00;
Memory[13386] = 8'h32;
Memory[13385] = 8'h22;
Memory[13384] = 8'hB3;
Memory[13391] = 8'h00;
Memory[13390] = 8'h02;
Memory[13389] = 8'h84;
Memory[13388] = 8'h63;
Memory[13395] = 8'h14;
Memory[13394] = 8'h00;
Memory[13393] = 8'h50;
Memory[13392] = 8'h6F;
Memory[13399] = 8'h22;
Memory[13398] = 8'h4C;
Memory[13397] = 8'hA2;
Memory[13396] = 8'h03;
Memory[13403] = 8'h00;
Memory[13402] = 8'h32;
Memory[13401] = 8'h22;
Memory[13400] = 8'hB3;
Memory[13407] = 8'h00;
Memory[13406] = 8'h02;
Memory[13405] = 8'h84;
Memory[13404] = 8'h63;
Memory[13411] = 8'h13;
Memory[13410] = 8'h40;
Memory[13409] = 8'h50;
Memory[13408] = 8'h6F;
Memory[13415] = 8'h22;
Memory[13414] = 8'h0C;
Memory[13413] = 8'hA2;
Memory[13412] = 8'h03;
Memory[13419] = 8'h00;
Memory[13418] = 8'h32;
Memory[13417] = 8'h22;
Memory[13416] = 8'hB3;
Memory[13423] = 8'h00;
Memory[13422] = 8'h02;
Memory[13421] = 8'h84;
Memory[13420] = 8'h63;
Memory[13427] = 8'h12;
Memory[13426] = 8'h80;
Memory[13425] = 8'h50;
Memory[13424] = 8'h6F;
Memory[13431] = 8'h21;
Memory[13430] = 8'hCC;
Memory[13429] = 8'hA2;
Memory[13428] = 8'h03;
Memory[13435] = 8'h00;
Memory[13434] = 8'h32;
Memory[13433] = 8'h22;
Memory[13432] = 8'hB3;
Memory[13439] = 8'h00;
Memory[13438] = 8'h02;
Memory[13437] = 8'h84;
Memory[13436] = 8'h63;
Memory[13443] = 8'h11;
Memory[13442] = 8'hC0;
Memory[13441] = 8'h50;
Memory[13440] = 8'h6F;
Memory[13447] = 8'h21;
Memory[13446] = 8'h8C;
Memory[13445] = 8'hA2;
Memory[13444] = 8'h03;
Memory[13451] = 8'h00;
Memory[13450] = 8'h32;
Memory[13449] = 8'h22;
Memory[13448] = 8'hB3;
Memory[13455] = 8'h00;
Memory[13454] = 8'h02;
Memory[13453] = 8'h84;
Memory[13452] = 8'h63;
Memory[13459] = 8'h11;
Memory[13458] = 8'h00;
Memory[13457] = 8'h50;
Memory[13456] = 8'h6F;
Memory[13463] = 8'h21;
Memory[13462] = 8'h4C;
Memory[13461] = 8'hA2;
Memory[13460] = 8'h03;
Memory[13467] = 8'h00;
Memory[13466] = 8'h32;
Memory[13465] = 8'h22;
Memory[13464] = 8'hB3;
Memory[13471] = 8'h00;
Memory[13470] = 8'h02;
Memory[13469] = 8'h84;
Memory[13468] = 8'h63;
Memory[13475] = 8'h10;
Memory[13474] = 8'h40;
Memory[13473] = 8'h50;
Memory[13472] = 8'h6F;
Memory[13479] = 8'h21;
Memory[13478] = 8'h0C;
Memory[13477] = 8'hA2;
Memory[13476] = 8'h03;
Memory[13483] = 8'h00;
Memory[13482] = 8'h32;
Memory[13481] = 8'h22;
Memory[13480] = 8'hB3;
Memory[13487] = 8'h00;
Memory[13486] = 8'h02;
Memory[13485] = 8'h84;
Memory[13484] = 8'h63;
Memory[13491] = 8'h0F;
Memory[13490] = 8'h80;
Memory[13489] = 8'h50;
Memory[13488] = 8'h6F;
Memory[13495] = 8'h20;
Memory[13494] = 8'hCC;
Memory[13493] = 8'hA2;
Memory[13492] = 8'h03;
Memory[13499] = 8'h00;
Memory[13498] = 8'h32;
Memory[13497] = 8'h22;
Memory[13496] = 8'hB3;
Memory[13503] = 8'h00;
Memory[13502] = 8'h02;
Memory[13501] = 8'h84;
Memory[13500] = 8'h63;
Memory[13507] = 8'h0E;
Memory[13506] = 8'hC0;
Memory[13505] = 8'h50;
Memory[13504] = 8'h6F;
Memory[13511] = 8'h20;
Memory[13510] = 8'h8C;
Memory[13509] = 8'hA2;
Memory[13508] = 8'h03;
Memory[13515] = 8'h00;
Memory[13514] = 8'h32;
Memory[13513] = 8'h22;
Memory[13512] = 8'hB3;
Memory[13519] = 8'h00;
Memory[13518] = 8'h02;
Memory[13517] = 8'h84;
Memory[13516] = 8'h63;
Memory[13523] = 8'h0E;
Memory[13522] = 8'h00;
Memory[13521] = 8'h50;
Memory[13520] = 8'h6F;
Memory[13527] = 8'h20;
Memory[13526] = 8'h4C;
Memory[13525] = 8'hA2;
Memory[13524] = 8'h03;
Memory[13531] = 8'h00;
Memory[13530] = 8'h32;
Memory[13529] = 8'h22;
Memory[13528] = 8'hB3;
Memory[13535] = 8'h00;
Memory[13534] = 8'h02;
Memory[13533] = 8'h84;
Memory[13532] = 8'h63;
Memory[13539] = 8'h0D;
Memory[13538] = 8'h40;
Memory[13537] = 8'h50;
Memory[13536] = 8'h6F;
Memory[13543] = 8'h20;
Memory[13542] = 8'h0C;
Memory[13541] = 8'hA2;
Memory[13540] = 8'h03;
Memory[13547] = 8'h00;
Memory[13546] = 8'h32;
Memory[13545] = 8'h22;
Memory[13544] = 8'hB3;
Memory[13551] = 8'h00;
Memory[13550] = 8'h02;
Memory[13549] = 8'h84;
Memory[13548] = 8'h63;
Memory[13555] = 8'h0C;
Memory[13554] = 8'h80;
Memory[13553] = 8'h50;
Memory[13552] = 8'h6F;
Memory[13559] = 8'h1F;
Memory[13558] = 8'hCC;
Memory[13557] = 8'hA2;
Memory[13556] = 8'h03;
Memory[13563] = 8'h00;
Memory[13562] = 8'h32;
Memory[13561] = 8'h22;
Memory[13560] = 8'hB3;
Memory[13567] = 8'h00;
Memory[13566] = 8'h02;
Memory[13565] = 8'h84;
Memory[13564] = 8'h63;
Memory[13571] = 8'h0B;
Memory[13570] = 8'hC0;
Memory[13569] = 8'h50;
Memory[13568] = 8'h6F;
Memory[13575] = 8'h1F;
Memory[13574] = 8'h8C;
Memory[13573] = 8'hA2;
Memory[13572] = 8'h03;
Memory[13579] = 8'h00;
Memory[13578] = 8'h32;
Memory[13577] = 8'h22;
Memory[13576] = 8'hB3;
Memory[13583] = 8'h00;
Memory[13582] = 8'h02;
Memory[13581] = 8'h84;
Memory[13580] = 8'h63;
Memory[13587] = 8'h0B;
Memory[13586] = 8'h00;
Memory[13585] = 8'h50;
Memory[13584] = 8'h6F;
Memory[13591] = 8'h1F;
Memory[13590] = 8'h4C;
Memory[13589] = 8'hA2;
Memory[13588] = 8'h03;
Memory[13595] = 8'h00;
Memory[13594] = 8'h32;
Memory[13593] = 8'h22;
Memory[13592] = 8'hB3;
Memory[13599] = 8'h00;
Memory[13598] = 8'h02;
Memory[13597] = 8'h84;
Memory[13596] = 8'h63;
Memory[13603] = 8'h0A;
Memory[13602] = 8'h40;
Memory[13601] = 8'h50;
Memory[13600] = 8'h6F;
Memory[13607] = 8'h1F;
Memory[13606] = 8'h0C;
Memory[13605] = 8'hA2;
Memory[13604] = 8'h03;
Memory[13611] = 8'h00;
Memory[13610] = 8'h32;
Memory[13609] = 8'h22;
Memory[13608] = 8'hB3;
Memory[13615] = 8'h00;
Memory[13614] = 8'h02;
Memory[13613] = 8'h84;
Memory[13612] = 8'h63;
Memory[13619] = 8'h09;
Memory[13618] = 8'h80;
Memory[13617] = 8'h50;
Memory[13616] = 8'h6F;
Memory[13623] = 8'h1E;
Memory[13622] = 8'hCC;
Memory[13621] = 8'hA2;
Memory[13620] = 8'h03;
Memory[13627] = 8'h00;
Memory[13626] = 8'h32;
Memory[13625] = 8'h22;
Memory[13624] = 8'hB3;
Memory[13631] = 8'h00;
Memory[13630] = 8'h02;
Memory[13629] = 8'h84;
Memory[13628] = 8'h63;
Memory[13635] = 8'h08;
Memory[13634] = 8'hC0;
Memory[13633] = 8'h50;
Memory[13632] = 8'h6F;
Memory[13639] = 8'h1E;
Memory[13638] = 8'h8C;
Memory[13637] = 8'hA2;
Memory[13636] = 8'h03;
Memory[13643] = 8'h00;
Memory[13642] = 8'h32;
Memory[13641] = 8'h22;
Memory[13640] = 8'hB3;
Memory[13647] = 8'h00;
Memory[13646] = 8'h02;
Memory[13645] = 8'h84;
Memory[13644] = 8'h63;
Memory[13651] = 8'h08;
Memory[13650] = 8'h00;
Memory[13649] = 8'h50;
Memory[13648] = 8'h6F;
Memory[13655] = 8'h1E;
Memory[13654] = 8'h4C;
Memory[13653] = 8'hA2;
Memory[13652] = 8'h03;
Memory[13659] = 8'h00;
Memory[13658] = 8'h32;
Memory[13657] = 8'h22;
Memory[13656] = 8'hB3;
Memory[13663] = 8'h00;
Memory[13662] = 8'h02;
Memory[13661] = 8'h84;
Memory[13660] = 8'h63;
Memory[13667] = 8'h07;
Memory[13666] = 8'h40;
Memory[13665] = 8'h50;
Memory[13664] = 8'h6F;
Memory[13671] = 8'h1E;
Memory[13670] = 8'h0C;
Memory[13669] = 8'hA2;
Memory[13668] = 8'h03;
Memory[13675] = 8'h00;
Memory[13674] = 8'h32;
Memory[13673] = 8'h22;
Memory[13672] = 8'hB3;
Memory[13679] = 8'h00;
Memory[13678] = 8'h02;
Memory[13677] = 8'h84;
Memory[13676] = 8'h63;
Memory[13683] = 8'h06;
Memory[13682] = 8'h80;
Memory[13681] = 8'h50;
Memory[13680] = 8'h6F;
Memory[13687] = 8'h1D;
Memory[13686] = 8'hCC;
Memory[13685] = 8'hA2;
Memory[13684] = 8'h03;
Memory[13691] = 8'h00;
Memory[13690] = 8'h32;
Memory[13689] = 8'h22;
Memory[13688] = 8'hB3;
Memory[13695] = 8'h00;
Memory[13694] = 8'h02;
Memory[13693] = 8'h84;
Memory[13692] = 8'h63;
Memory[13699] = 8'h05;
Memory[13698] = 8'hC0;
Memory[13697] = 8'h50;
Memory[13696] = 8'h6F;
Memory[13703] = 8'h1D;
Memory[13702] = 8'h8C;
Memory[13701] = 8'hA2;
Memory[13700] = 8'h03;
Memory[13707] = 8'h00;
Memory[13706] = 8'h32;
Memory[13705] = 8'h22;
Memory[13704] = 8'hB3;
Memory[13711] = 8'h00;
Memory[13710] = 8'h02;
Memory[13709] = 8'h84;
Memory[13708] = 8'h63;
Memory[13715] = 8'h05;
Memory[13714] = 8'h00;
Memory[13713] = 8'h50;
Memory[13712] = 8'h6F;
Memory[13719] = 8'h1D;
Memory[13718] = 8'h4C;
Memory[13717] = 8'hA2;
Memory[13716] = 8'h03;
Memory[13723] = 8'h00;
Memory[13722] = 8'h32;
Memory[13721] = 8'h22;
Memory[13720] = 8'hB3;
Memory[13727] = 8'h00;
Memory[13726] = 8'h02;
Memory[13725] = 8'h84;
Memory[13724] = 8'h63;
Memory[13731] = 8'h04;
Memory[13730] = 8'h40;
Memory[13729] = 8'h50;
Memory[13728] = 8'h6F;
Memory[13735] = 8'h1D;
Memory[13734] = 8'h0C;
Memory[13733] = 8'hA2;
Memory[13732] = 8'h03;
Memory[13739] = 8'h00;
Memory[13738] = 8'h32;
Memory[13737] = 8'h22;
Memory[13736] = 8'hB3;
Memory[13743] = 8'h00;
Memory[13742] = 8'h02;
Memory[13741] = 8'h84;
Memory[13740] = 8'h63;
Memory[13747] = 8'h03;
Memory[13746] = 8'h80;
Memory[13745] = 8'h50;
Memory[13744] = 8'h6F;
Memory[13751] = 8'h1C;
Memory[13750] = 8'hCC;
Memory[13749] = 8'hA2;
Memory[13748] = 8'h03;
Memory[13755] = 8'h00;
Memory[13754] = 8'h32;
Memory[13753] = 8'h22;
Memory[13752] = 8'hB3;
Memory[13759] = 8'h00;
Memory[13758] = 8'h02;
Memory[13757] = 8'h84;
Memory[13756] = 8'h63;
Memory[13763] = 8'h02;
Memory[13762] = 8'hC0;
Memory[13761] = 8'h50;
Memory[13760] = 8'h6F;
Memory[13767] = 8'h1C;
Memory[13766] = 8'h8C;
Memory[13765] = 8'hA2;
Memory[13764] = 8'h03;
Memory[13771] = 8'h00;
Memory[13770] = 8'h32;
Memory[13769] = 8'h22;
Memory[13768] = 8'hB3;
Memory[13775] = 8'h00;
Memory[13774] = 8'h02;
Memory[13773] = 8'h84;
Memory[13772] = 8'h63;
Memory[13779] = 8'h02;
Memory[13778] = 8'h00;
Memory[13777] = 8'h50;
Memory[13776] = 8'h6F;
Memory[13783] = 8'h1C;
Memory[13782] = 8'h4C;
Memory[13781] = 8'hA2;
Memory[13780] = 8'h03;
Memory[13787] = 8'h00;
Memory[13786] = 8'h32;
Memory[13785] = 8'h22;
Memory[13784] = 8'hB3;
Memory[13791] = 8'h00;
Memory[13790] = 8'h02;
Memory[13789] = 8'h84;
Memory[13788] = 8'h63;
Memory[13795] = 8'h01;
Memory[13794] = 8'h40;
Memory[13793] = 8'h50;
Memory[13792] = 8'h6F;
Memory[13799] = 8'h1C;
Memory[13798] = 8'h0C;
Memory[13797] = 8'hA2;
Memory[13796] = 8'h03;
Memory[13803] = 8'h00;
Memory[13802] = 8'h32;
Memory[13801] = 8'h22;
Memory[13800] = 8'hB3;
Memory[13807] = 8'h00;
Memory[13806] = 8'h02;
Memory[13805] = 8'h84;
Memory[13804] = 8'h63;
Memory[13811] = 8'h00;
Memory[13810] = 8'h80;
Memory[13809] = 8'h50;
Memory[13808] = 8'h6F;
Memory[13815] = 8'h1B;
Memory[13814] = 8'hCC;
Memory[13813] = 8'hA2;
Memory[13812] = 8'h03;
Memory[13819] = 8'h00;
Memory[13818] = 8'h32;
Memory[13817] = 8'h22;
Memory[13816] = 8'hB3;
Memory[13823] = 8'h00;
Memory[13822] = 8'h02;
Memory[13821] = 8'h84;
Memory[13820] = 8'h63;
Memory[13827] = 8'h7F;
Memory[13826] = 8'hD0;
Memory[13825] = 8'h40;
Memory[13824] = 8'h6F;
Memory[13831] = 8'h1B;
Memory[13830] = 8'h8C;
Memory[13829] = 8'hA2;
Memory[13828] = 8'h03;
Memory[13835] = 8'h00;
Memory[13834] = 8'h32;
Memory[13833] = 8'h22;
Memory[13832] = 8'hB3;
Memory[13839] = 8'h00;
Memory[13838] = 8'h02;
Memory[13837] = 8'h84;
Memory[13836] = 8'h63;
Memory[13843] = 8'h7F;
Memory[13842] = 8'h10;
Memory[13841] = 8'h40;
Memory[13840] = 8'h6F;
Memory[13847] = 8'h1B;
Memory[13846] = 8'h4C;
Memory[13845] = 8'hA2;
Memory[13844] = 8'h03;
Memory[13851] = 8'h00;
Memory[13850] = 8'h32;
Memory[13849] = 8'h22;
Memory[13848] = 8'hB3;
Memory[13855] = 8'h00;
Memory[13854] = 8'h02;
Memory[13853] = 8'h84;
Memory[13852] = 8'h63;
Memory[13859] = 8'h7E;
Memory[13858] = 8'h50;
Memory[13857] = 8'h40;
Memory[13856] = 8'h6F;
Memory[13863] = 8'h1B;
Memory[13862] = 8'h0C;
Memory[13861] = 8'hA2;
Memory[13860] = 8'h03;
Memory[13867] = 8'h00;
Memory[13866] = 8'h32;
Memory[13865] = 8'h22;
Memory[13864] = 8'hB3;
Memory[13871] = 8'h00;
Memory[13870] = 8'h02;
Memory[13869] = 8'h84;
Memory[13868] = 8'h63;
Memory[13875] = 8'h7D;
Memory[13874] = 8'h90;
Memory[13873] = 8'h40;
Memory[13872] = 8'h6F;
Memory[13879] = 8'h1A;
Memory[13878] = 8'hCC;
Memory[13877] = 8'hA2;
Memory[13876] = 8'h03;
Memory[13883] = 8'h00;
Memory[13882] = 8'h32;
Memory[13881] = 8'h22;
Memory[13880] = 8'hB3;
Memory[13887] = 8'h00;
Memory[13886] = 8'h02;
Memory[13885] = 8'h84;
Memory[13884] = 8'h63;
Memory[13891] = 8'h7C;
Memory[13890] = 8'hD0;
Memory[13889] = 8'h40;
Memory[13888] = 8'h6F;
Memory[13895] = 8'h1A;
Memory[13894] = 8'h8C;
Memory[13893] = 8'hA2;
Memory[13892] = 8'h03;
Memory[13899] = 8'h00;
Memory[13898] = 8'h32;
Memory[13897] = 8'h22;
Memory[13896] = 8'hB3;
Memory[13903] = 8'h00;
Memory[13902] = 8'h02;
Memory[13901] = 8'h84;
Memory[13900] = 8'h63;
Memory[13907] = 8'h7C;
Memory[13906] = 8'h10;
Memory[13905] = 8'h40;
Memory[13904] = 8'h6F;
Memory[13911] = 8'h1A;
Memory[13910] = 8'h4C;
Memory[13909] = 8'hA2;
Memory[13908] = 8'h03;
Memory[13915] = 8'h00;
Memory[13914] = 8'h32;
Memory[13913] = 8'h22;
Memory[13912] = 8'hB3;
Memory[13919] = 8'h00;
Memory[13918] = 8'h02;
Memory[13917] = 8'h84;
Memory[13916] = 8'h63;
Memory[13923] = 8'h7B;
Memory[13922] = 8'h50;
Memory[13921] = 8'h40;
Memory[13920] = 8'h6F;
Memory[13927] = 8'h1A;
Memory[13926] = 8'h0C;
Memory[13925] = 8'hA2;
Memory[13924] = 8'h03;
Memory[13931] = 8'h00;
Memory[13930] = 8'h32;
Memory[13929] = 8'h22;
Memory[13928] = 8'hB3;
Memory[13935] = 8'h00;
Memory[13934] = 8'h02;
Memory[13933] = 8'h84;
Memory[13932] = 8'h63;
Memory[13939] = 8'h7A;
Memory[13938] = 8'h90;
Memory[13937] = 8'h40;
Memory[13936] = 8'h6F;
Memory[13943] = 8'h19;
Memory[13942] = 8'hCC;
Memory[13941] = 8'hA2;
Memory[13940] = 8'h03;
Memory[13947] = 8'h00;
Memory[13946] = 8'h32;
Memory[13945] = 8'h22;
Memory[13944] = 8'hB3;
Memory[13951] = 8'h00;
Memory[13950] = 8'h02;
Memory[13949] = 8'h84;
Memory[13948] = 8'h63;
Memory[13955] = 8'h79;
Memory[13954] = 8'hD0;
Memory[13953] = 8'h40;
Memory[13952] = 8'h6F;
Memory[13959] = 8'h19;
Memory[13958] = 8'h8C;
Memory[13957] = 8'hA2;
Memory[13956] = 8'h03;
Memory[13963] = 8'h00;
Memory[13962] = 8'h32;
Memory[13961] = 8'h22;
Memory[13960] = 8'hB3;
Memory[13967] = 8'h00;
Memory[13966] = 8'h02;
Memory[13965] = 8'h84;
Memory[13964] = 8'h63;
Memory[13971] = 8'h79;
Memory[13970] = 8'h10;
Memory[13969] = 8'h40;
Memory[13968] = 8'h6F;
Memory[13975] = 8'h19;
Memory[13974] = 8'h4C;
Memory[13973] = 8'hA2;
Memory[13972] = 8'h03;
Memory[13979] = 8'h00;
Memory[13978] = 8'h32;
Memory[13977] = 8'h22;
Memory[13976] = 8'hB3;
Memory[13983] = 8'h00;
Memory[13982] = 8'h02;
Memory[13981] = 8'h84;
Memory[13980] = 8'h63;
Memory[13987] = 8'h78;
Memory[13986] = 8'h50;
Memory[13985] = 8'h40;
Memory[13984] = 8'h6F;
Memory[13991] = 8'h19;
Memory[13990] = 8'h0C;
Memory[13989] = 8'hA2;
Memory[13988] = 8'h03;
Memory[13995] = 8'h00;
Memory[13994] = 8'h32;
Memory[13993] = 8'h22;
Memory[13992] = 8'hB3;
Memory[13999] = 8'h00;
Memory[13998] = 8'h02;
Memory[13997] = 8'h84;
Memory[13996] = 8'h63;
Memory[14003] = 8'h77;
Memory[14002] = 8'h90;
Memory[14001] = 8'h40;
Memory[14000] = 8'h6F;
Memory[14007] = 8'h18;
Memory[14006] = 8'hCC;
Memory[14005] = 8'hA2;
Memory[14004] = 8'h03;
Memory[14011] = 8'h00;
Memory[14010] = 8'h32;
Memory[14009] = 8'h22;
Memory[14008] = 8'hB3;
Memory[14015] = 8'h00;
Memory[14014] = 8'h02;
Memory[14013] = 8'h84;
Memory[14012] = 8'h63;
Memory[14019] = 8'h76;
Memory[14018] = 8'hD0;
Memory[14017] = 8'h40;
Memory[14016] = 8'h6F;
Memory[14023] = 8'h18;
Memory[14022] = 8'h8C;
Memory[14021] = 8'hA2;
Memory[14020] = 8'h03;
Memory[14027] = 8'h00;
Memory[14026] = 8'h32;
Memory[14025] = 8'h22;
Memory[14024] = 8'hB3;
Memory[14031] = 8'h00;
Memory[14030] = 8'h02;
Memory[14029] = 8'h84;
Memory[14028] = 8'h63;
Memory[14035] = 8'h76;
Memory[14034] = 8'h10;
Memory[14033] = 8'h40;
Memory[14032] = 8'h6F;
Memory[14039] = 8'h18;
Memory[14038] = 8'h4C;
Memory[14037] = 8'hA2;
Memory[14036] = 8'h03;
Memory[14043] = 8'h00;
Memory[14042] = 8'h32;
Memory[14041] = 8'h22;
Memory[14040] = 8'hB3;
Memory[14047] = 8'h00;
Memory[14046] = 8'h02;
Memory[14045] = 8'h84;
Memory[14044] = 8'h63;
Memory[14051] = 8'h75;
Memory[14050] = 8'h50;
Memory[14049] = 8'h40;
Memory[14048] = 8'h6F;
Memory[14055] = 8'h18;
Memory[14054] = 8'h0C;
Memory[14053] = 8'hA2;
Memory[14052] = 8'h03;
Memory[14059] = 8'h00;
Memory[14058] = 8'h32;
Memory[14057] = 8'h22;
Memory[14056] = 8'hB3;
Memory[14063] = 8'h00;
Memory[14062] = 8'h02;
Memory[14061] = 8'h84;
Memory[14060] = 8'h63;
Memory[14067] = 8'h74;
Memory[14066] = 8'h90;
Memory[14065] = 8'h40;
Memory[14064] = 8'h6F;
Memory[14071] = 8'h17;
Memory[14070] = 8'hCC;
Memory[14069] = 8'hA2;
Memory[14068] = 8'h03;
Memory[14075] = 8'h00;
Memory[14074] = 8'h32;
Memory[14073] = 8'h22;
Memory[14072] = 8'hB3;
Memory[14079] = 8'h00;
Memory[14078] = 8'h02;
Memory[14077] = 8'h84;
Memory[14076] = 8'h63;
Memory[14083] = 8'h73;
Memory[14082] = 8'hD0;
Memory[14081] = 8'h40;
Memory[14080] = 8'h6F;
Memory[14087] = 8'h17;
Memory[14086] = 8'h8C;
Memory[14085] = 8'hA2;
Memory[14084] = 8'h03;
Memory[14091] = 8'h00;
Memory[14090] = 8'h32;
Memory[14089] = 8'h22;
Memory[14088] = 8'hB3;
Memory[14095] = 8'h00;
Memory[14094] = 8'h02;
Memory[14093] = 8'h84;
Memory[14092] = 8'h63;
Memory[14099] = 8'h73;
Memory[14098] = 8'h10;
Memory[14097] = 8'h40;
Memory[14096] = 8'h6F;
Memory[14103] = 8'h17;
Memory[14102] = 8'h4C;
Memory[14101] = 8'hA2;
Memory[14100] = 8'h03;
Memory[14107] = 8'h00;
Memory[14106] = 8'h32;
Memory[14105] = 8'h22;
Memory[14104] = 8'hB3;
Memory[14111] = 8'h00;
Memory[14110] = 8'h02;
Memory[14109] = 8'h84;
Memory[14108] = 8'h63;
Memory[14115] = 8'h72;
Memory[14114] = 8'h50;
Memory[14113] = 8'h40;
Memory[14112] = 8'h6F;
Memory[14119] = 8'h17;
Memory[14118] = 8'h0C;
Memory[14117] = 8'hA2;
Memory[14116] = 8'h03;
Memory[14123] = 8'h00;
Memory[14122] = 8'h32;
Memory[14121] = 8'h22;
Memory[14120] = 8'hB3;
Memory[14127] = 8'h00;
Memory[14126] = 8'h02;
Memory[14125] = 8'h84;
Memory[14124] = 8'h63;
Memory[14131] = 8'h71;
Memory[14130] = 8'h90;
Memory[14129] = 8'h40;
Memory[14128] = 8'h6F;
Memory[14135] = 8'h16;
Memory[14134] = 8'hCC;
Memory[14133] = 8'hA2;
Memory[14132] = 8'h03;
Memory[14139] = 8'h00;
Memory[14138] = 8'h32;
Memory[14137] = 8'h22;
Memory[14136] = 8'hB3;
Memory[14143] = 8'h00;
Memory[14142] = 8'h02;
Memory[14141] = 8'h84;
Memory[14140] = 8'h63;
Memory[14147] = 8'h70;
Memory[14146] = 8'hD0;
Memory[14145] = 8'h40;
Memory[14144] = 8'h6F;
Memory[14151] = 8'h16;
Memory[14150] = 8'h8C;
Memory[14149] = 8'hA2;
Memory[14148] = 8'h03;
Memory[14155] = 8'h00;
Memory[14154] = 8'h32;
Memory[14153] = 8'h22;
Memory[14152] = 8'hB3;
Memory[14159] = 8'h00;
Memory[14158] = 8'h02;
Memory[14157] = 8'h84;
Memory[14156] = 8'h63;
Memory[14163] = 8'h70;
Memory[14162] = 8'h10;
Memory[14161] = 8'h40;
Memory[14160] = 8'h6F;
Memory[14167] = 8'h16;
Memory[14166] = 8'h4C;
Memory[14165] = 8'hA2;
Memory[14164] = 8'h03;
Memory[14171] = 8'h00;
Memory[14170] = 8'h32;
Memory[14169] = 8'h22;
Memory[14168] = 8'hB3;
Memory[14175] = 8'h00;
Memory[14174] = 8'h02;
Memory[14173] = 8'h84;
Memory[14172] = 8'h63;
Memory[14179] = 8'h6F;
Memory[14178] = 8'h50;
Memory[14177] = 8'h40;
Memory[14176] = 8'h6F;
Memory[14183] = 8'h16;
Memory[14182] = 8'h0C;
Memory[14181] = 8'hA2;
Memory[14180] = 8'h03;
Memory[14187] = 8'h00;
Memory[14186] = 8'h32;
Memory[14185] = 8'h22;
Memory[14184] = 8'hB3;
Memory[14191] = 8'h00;
Memory[14190] = 8'h02;
Memory[14189] = 8'h84;
Memory[14188] = 8'h63;
Memory[14195] = 8'h6E;
Memory[14194] = 8'h90;
Memory[14193] = 8'h40;
Memory[14192] = 8'h6F;
Memory[14199] = 8'h15;
Memory[14198] = 8'hCC;
Memory[14197] = 8'hA2;
Memory[14196] = 8'h03;
Memory[14203] = 8'h00;
Memory[14202] = 8'h32;
Memory[14201] = 8'h22;
Memory[14200] = 8'hB3;
Memory[14207] = 8'h00;
Memory[14206] = 8'h02;
Memory[14205] = 8'h84;
Memory[14204] = 8'h63;
Memory[14211] = 8'h6D;
Memory[14210] = 8'hD0;
Memory[14209] = 8'h40;
Memory[14208] = 8'h6F;
Memory[14215] = 8'h15;
Memory[14214] = 8'h8C;
Memory[14213] = 8'hA2;
Memory[14212] = 8'h03;
Memory[14219] = 8'h00;
Memory[14218] = 8'h32;
Memory[14217] = 8'h22;
Memory[14216] = 8'hB3;
Memory[14223] = 8'h00;
Memory[14222] = 8'h02;
Memory[14221] = 8'h84;
Memory[14220] = 8'h63;
Memory[14227] = 8'h6D;
Memory[14226] = 8'h10;
Memory[14225] = 8'h40;
Memory[14224] = 8'h6F;
Memory[14231] = 8'h15;
Memory[14230] = 8'h4C;
Memory[14229] = 8'hA2;
Memory[14228] = 8'h03;
Memory[14235] = 8'h00;
Memory[14234] = 8'h32;
Memory[14233] = 8'h22;
Memory[14232] = 8'hB3;
Memory[14239] = 8'h00;
Memory[14238] = 8'h02;
Memory[14237] = 8'h84;
Memory[14236] = 8'h63;
Memory[14243] = 8'h6C;
Memory[14242] = 8'h50;
Memory[14241] = 8'h40;
Memory[14240] = 8'h6F;
Memory[14247] = 8'h15;
Memory[14246] = 8'h0C;
Memory[14245] = 8'hA2;
Memory[14244] = 8'h03;
Memory[14251] = 8'h00;
Memory[14250] = 8'h32;
Memory[14249] = 8'h22;
Memory[14248] = 8'hB3;
Memory[14255] = 8'h00;
Memory[14254] = 8'h02;
Memory[14253] = 8'h84;
Memory[14252] = 8'h63;
Memory[14259] = 8'h6B;
Memory[14258] = 8'h90;
Memory[14257] = 8'h40;
Memory[14256] = 8'h6F;
Memory[14263] = 8'h14;
Memory[14262] = 8'hCC;
Memory[14261] = 8'hA2;
Memory[14260] = 8'h03;
Memory[14267] = 8'h00;
Memory[14266] = 8'h32;
Memory[14265] = 8'h22;
Memory[14264] = 8'hB3;
Memory[14271] = 8'h00;
Memory[14270] = 8'h02;
Memory[14269] = 8'h84;
Memory[14268] = 8'h63;
Memory[14275] = 8'h6A;
Memory[14274] = 8'hD0;
Memory[14273] = 8'h40;
Memory[14272] = 8'h6F;
Memory[14279] = 8'h14;
Memory[14278] = 8'h8C;
Memory[14277] = 8'hA2;
Memory[14276] = 8'h03;
Memory[14283] = 8'h00;
Memory[14282] = 8'h32;
Memory[14281] = 8'h22;
Memory[14280] = 8'hB3;
Memory[14287] = 8'h00;
Memory[14286] = 8'h02;
Memory[14285] = 8'h84;
Memory[14284] = 8'h63;
Memory[14291] = 8'h6A;
Memory[14290] = 8'h10;
Memory[14289] = 8'h40;
Memory[14288] = 8'h6F;
Memory[14295] = 8'h14;
Memory[14294] = 8'h4C;
Memory[14293] = 8'hA2;
Memory[14292] = 8'h03;
Memory[14299] = 8'h00;
Memory[14298] = 8'h32;
Memory[14297] = 8'h22;
Memory[14296] = 8'hB3;
Memory[14303] = 8'h00;
Memory[14302] = 8'h02;
Memory[14301] = 8'h84;
Memory[14300] = 8'h63;
Memory[14307] = 8'h69;
Memory[14306] = 8'h50;
Memory[14305] = 8'h40;
Memory[14304] = 8'h6F;
Memory[14311] = 8'h14;
Memory[14310] = 8'h0C;
Memory[14309] = 8'hA2;
Memory[14308] = 8'h03;
Memory[14315] = 8'h00;
Memory[14314] = 8'h32;
Memory[14313] = 8'h22;
Memory[14312] = 8'hB3;
Memory[14319] = 8'h00;
Memory[14318] = 8'h02;
Memory[14317] = 8'h84;
Memory[14316] = 8'h63;
Memory[14323] = 8'h68;
Memory[14322] = 8'h90;
Memory[14321] = 8'h40;
Memory[14320] = 8'h6F;
Memory[14327] = 8'h13;
Memory[14326] = 8'hCC;
Memory[14325] = 8'hA2;
Memory[14324] = 8'h03;
Memory[14331] = 8'h00;
Memory[14330] = 8'h32;
Memory[14329] = 8'h22;
Memory[14328] = 8'hB3;
Memory[14335] = 8'h00;
Memory[14334] = 8'h02;
Memory[14333] = 8'h84;
Memory[14332] = 8'h63;
Memory[14339] = 8'h67;
Memory[14338] = 8'hD0;
Memory[14337] = 8'h40;
Memory[14336] = 8'h6F;
Memory[14343] = 8'h13;
Memory[14342] = 8'h8C;
Memory[14341] = 8'hA2;
Memory[14340] = 8'h03;
Memory[14347] = 8'h00;
Memory[14346] = 8'h32;
Memory[14345] = 8'h22;
Memory[14344] = 8'hB3;
Memory[14351] = 8'h00;
Memory[14350] = 8'h02;
Memory[14349] = 8'h84;
Memory[14348] = 8'h63;
Memory[14355] = 8'h67;
Memory[14354] = 8'h10;
Memory[14353] = 8'h40;
Memory[14352] = 8'h6F;
Memory[14359] = 8'h13;
Memory[14358] = 8'h4C;
Memory[14357] = 8'hA2;
Memory[14356] = 8'h03;
Memory[14363] = 8'h00;
Memory[14362] = 8'h32;
Memory[14361] = 8'h22;
Memory[14360] = 8'hB3;
Memory[14367] = 8'h00;
Memory[14366] = 8'h02;
Memory[14365] = 8'h84;
Memory[14364] = 8'h63;
Memory[14371] = 8'h66;
Memory[14370] = 8'h50;
Memory[14369] = 8'h40;
Memory[14368] = 8'h6F;
Memory[14375] = 8'h13;
Memory[14374] = 8'h0C;
Memory[14373] = 8'hA2;
Memory[14372] = 8'h03;
Memory[14379] = 8'h00;
Memory[14378] = 8'h32;
Memory[14377] = 8'h22;
Memory[14376] = 8'hB3;
Memory[14383] = 8'h00;
Memory[14382] = 8'h02;
Memory[14381] = 8'h84;
Memory[14380] = 8'h63;
Memory[14387] = 8'h65;
Memory[14386] = 8'h90;
Memory[14385] = 8'h40;
Memory[14384] = 8'h6F;
Memory[14391] = 8'h12;
Memory[14390] = 8'hCC;
Memory[14389] = 8'hA2;
Memory[14388] = 8'h03;
Memory[14395] = 8'h00;
Memory[14394] = 8'h32;
Memory[14393] = 8'h22;
Memory[14392] = 8'hB3;
Memory[14399] = 8'h00;
Memory[14398] = 8'h02;
Memory[14397] = 8'h84;
Memory[14396] = 8'h63;
Memory[14403] = 8'h64;
Memory[14402] = 8'hD0;
Memory[14401] = 8'h40;
Memory[14400] = 8'h6F;
Memory[14407] = 8'h12;
Memory[14406] = 8'h8C;
Memory[14405] = 8'hA2;
Memory[14404] = 8'h03;
Memory[14411] = 8'h00;
Memory[14410] = 8'h32;
Memory[14409] = 8'h22;
Memory[14408] = 8'hB3;
Memory[14415] = 8'h00;
Memory[14414] = 8'h02;
Memory[14413] = 8'h84;
Memory[14412] = 8'h63;
Memory[14419] = 8'h64;
Memory[14418] = 8'h10;
Memory[14417] = 8'h40;
Memory[14416] = 8'h6F;
Memory[14423] = 8'h12;
Memory[14422] = 8'h4C;
Memory[14421] = 8'hA2;
Memory[14420] = 8'h03;
Memory[14427] = 8'h00;
Memory[14426] = 8'h32;
Memory[14425] = 8'h22;
Memory[14424] = 8'hB3;
Memory[14431] = 8'h00;
Memory[14430] = 8'h02;
Memory[14429] = 8'h84;
Memory[14428] = 8'h63;
Memory[14435] = 8'h63;
Memory[14434] = 8'h50;
Memory[14433] = 8'h40;
Memory[14432] = 8'h6F;
Memory[14439] = 8'h12;
Memory[14438] = 8'h0C;
Memory[14437] = 8'hA2;
Memory[14436] = 8'h03;
Memory[14443] = 8'h00;
Memory[14442] = 8'h32;
Memory[14441] = 8'h22;
Memory[14440] = 8'hB3;
Memory[14447] = 8'h00;
Memory[14446] = 8'h02;
Memory[14445] = 8'h84;
Memory[14444] = 8'h63;
Memory[14451] = 8'h62;
Memory[14450] = 8'h90;
Memory[14449] = 8'h40;
Memory[14448] = 8'h6F;
Memory[14455] = 8'h11;
Memory[14454] = 8'hCC;
Memory[14453] = 8'hA2;
Memory[14452] = 8'h03;
Memory[14459] = 8'h00;
Memory[14458] = 8'h32;
Memory[14457] = 8'h22;
Memory[14456] = 8'hB3;
Memory[14463] = 8'h00;
Memory[14462] = 8'h02;
Memory[14461] = 8'h84;
Memory[14460] = 8'h63;
Memory[14467] = 8'h61;
Memory[14466] = 8'hD0;
Memory[14465] = 8'h40;
Memory[14464] = 8'h6F;
Memory[14471] = 8'h11;
Memory[14470] = 8'h8C;
Memory[14469] = 8'hA2;
Memory[14468] = 8'h03;
Memory[14475] = 8'h00;
Memory[14474] = 8'h32;
Memory[14473] = 8'h22;
Memory[14472] = 8'hB3;
Memory[14479] = 8'h00;
Memory[14478] = 8'h02;
Memory[14477] = 8'h84;
Memory[14476] = 8'h63;
Memory[14483] = 8'h61;
Memory[14482] = 8'h10;
Memory[14481] = 8'h40;
Memory[14480] = 8'h6F;
Memory[14487] = 8'h11;
Memory[14486] = 8'h4C;
Memory[14485] = 8'hA2;
Memory[14484] = 8'h03;
Memory[14491] = 8'h00;
Memory[14490] = 8'h32;
Memory[14489] = 8'h22;
Memory[14488] = 8'hB3;
Memory[14495] = 8'h00;
Memory[14494] = 8'h02;
Memory[14493] = 8'h84;
Memory[14492] = 8'h63;
Memory[14499] = 8'h60;
Memory[14498] = 8'h50;
Memory[14497] = 8'h40;
Memory[14496] = 8'h6F;
Memory[14503] = 8'h11;
Memory[14502] = 8'h0C;
Memory[14501] = 8'hA2;
Memory[14500] = 8'h03;
Memory[14507] = 8'h00;
Memory[14506] = 8'h32;
Memory[14505] = 8'h22;
Memory[14504] = 8'hB3;
Memory[14511] = 8'h00;
Memory[14510] = 8'h02;
Memory[14509] = 8'h84;
Memory[14508] = 8'h63;
Memory[14515] = 8'h5F;
Memory[14514] = 8'h90;
Memory[14513] = 8'h40;
Memory[14512] = 8'h6F;
Memory[14519] = 8'h10;
Memory[14518] = 8'hCC;
Memory[14517] = 8'hA2;
Memory[14516] = 8'h03;
Memory[14523] = 8'h00;
Memory[14522] = 8'h32;
Memory[14521] = 8'h22;
Memory[14520] = 8'hB3;
Memory[14527] = 8'h00;
Memory[14526] = 8'h02;
Memory[14525] = 8'h84;
Memory[14524] = 8'h63;
Memory[14531] = 8'h5E;
Memory[14530] = 8'hD0;
Memory[14529] = 8'h40;
Memory[14528] = 8'h6F;
Memory[14535] = 8'h10;
Memory[14534] = 8'h8C;
Memory[14533] = 8'hA2;
Memory[14532] = 8'h03;
Memory[14539] = 8'h00;
Memory[14538] = 8'h32;
Memory[14537] = 8'h22;
Memory[14536] = 8'hB3;
Memory[14543] = 8'h00;
Memory[14542] = 8'h02;
Memory[14541] = 8'h84;
Memory[14540] = 8'h63;
Memory[14547] = 8'h5E;
Memory[14546] = 8'h10;
Memory[14545] = 8'h40;
Memory[14544] = 8'h6F;
Memory[14551] = 8'h10;
Memory[14550] = 8'h4C;
Memory[14549] = 8'hA2;
Memory[14548] = 8'h03;
Memory[14555] = 8'h00;
Memory[14554] = 8'h32;
Memory[14553] = 8'h22;
Memory[14552] = 8'hB3;
Memory[14559] = 8'h00;
Memory[14558] = 8'h02;
Memory[14557] = 8'h84;
Memory[14556] = 8'h63;
Memory[14563] = 8'h5D;
Memory[14562] = 8'h50;
Memory[14561] = 8'h40;
Memory[14560] = 8'h6F;
Memory[14567] = 8'h10;
Memory[14566] = 8'h0C;
Memory[14565] = 8'hA2;
Memory[14564] = 8'h03;
Memory[14571] = 8'h00;
Memory[14570] = 8'h32;
Memory[14569] = 8'h22;
Memory[14568] = 8'hB3;
Memory[14575] = 8'h00;
Memory[14574] = 8'h02;
Memory[14573] = 8'h84;
Memory[14572] = 8'h63;
Memory[14579] = 8'h5C;
Memory[14578] = 8'h90;
Memory[14577] = 8'h40;
Memory[14576] = 8'h6F;
Memory[14583] = 8'h0F;
Memory[14582] = 8'hCC;
Memory[14581] = 8'hA2;
Memory[14580] = 8'h03;
Memory[14587] = 8'h00;
Memory[14586] = 8'h32;
Memory[14585] = 8'h22;
Memory[14584] = 8'hB3;
Memory[14591] = 8'h00;
Memory[14590] = 8'h02;
Memory[14589] = 8'h84;
Memory[14588] = 8'h63;
Memory[14595] = 8'h5B;
Memory[14594] = 8'hD0;
Memory[14593] = 8'h40;
Memory[14592] = 8'h6F;
Memory[14599] = 8'h0F;
Memory[14598] = 8'h8C;
Memory[14597] = 8'hA2;
Memory[14596] = 8'h03;
Memory[14603] = 8'h00;
Memory[14602] = 8'h32;
Memory[14601] = 8'h22;
Memory[14600] = 8'hB3;
Memory[14607] = 8'h00;
Memory[14606] = 8'h02;
Memory[14605] = 8'h84;
Memory[14604] = 8'h63;
Memory[14611] = 8'h5B;
Memory[14610] = 8'h10;
Memory[14609] = 8'h40;
Memory[14608] = 8'h6F;
Memory[14615] = 8'h0F;
Memory[14614] = 8'h4C;
Memory[14613] = 8'hA2;
Memory[14612] = 8'h03;
Memory[14619] = 8'h00;
Memory[14618] = 8'h32;
Memory[14617] = 8'h22;
Memory[14616] = 8'hB3;
Memory[14623] = 8'h00;
Memory[14622] = 8'h02;
Memory[14621] = 8'h84;
Memory[14620] = 8'h63;
Memory[14627] = 8'h5A;
Memory[14626] = 8'h50;
Memory[14625] = 8'h40;
Memory[14624] = 8'h6F;
Memory[14631] = 8'h0F;
Memory[14630] = 8'h0C;
Memory[14629] = 8'hA2;
Memory[14628] = 8'h03;
Memory[14635] = 8'h00;
Memory[14634] = 8'h32;
Memory[14633] = 8'h22;
Memory[14632] = 8'hB3;
Memory[14639] = 8'h00;
Memory[14638] = 8'h02;
Memory[14637] = 8'h84;
Memory[14636] = 8'h63;
Memory[14643] = 8'h59;
Memory[14642] = 8'h90;
Memory[14641] = 8'h40;
Memory[14640] = 8'h6F;
Memory[14647] = 8'h0E;
Memory[14646] = 8'hCC;
Memory[14645] = 8'hA2;
Memory[14644] = 8'h03;
Memory[14651] = 8'h00;
Memory[14650] = 8'h32;
Memory[14649] = 8'h22;
Memory[14648] = 8'hB3;
Memory[14655] = 8'h00;
Memory[14654] = 8'h02;
Memory[14653] = 8'h84;
Memory[14652] = 8'h63;
Memory[14659] = 8'h58;
Memory[14658] = 8'hD0;
Memory[14657] = 8'h40;
Memory[14656] = 8'h6F;
Memory[14663] = 8'h0E;
Memory[14662] = 8'h8C;
Memory[14661] = 8'hA2;
Memory[14660] = 8'h03;
Memory[14667] = 8'h00;
Memory[14666] = 8'h32;
Memory[14665] = 8'h22;
Memory[14664] = 8'hB3;
Memory[14671] = 8'h00;
Memory[14670] = 8'h02;
Memory[14669] = 8'h84;
Memory[14668] = 8'h63;
Memory[14675] = 8'h58;
Memory[14674] = 8'h10;
Memory[14673] = 8'h40;
Memory[14672] = 8'h6F;
Memory[14679] = 8'h0E;
Memory[14678] = 8'h4C;
Memory[14677] = 8'hA2;
Memory[14676] = 8'h03;
Memory[14683] = 8'h00;
Memory[14682] = 8'h32;
Memory[14681] = 8'h22;
Memory[14680] = 8'hB3;
Memory[14687] = 8'h00;
Memory[14686] = 8'h02;
Memory[14685] = 8'h84;
Memory[14684] = 8'h63;
Memory[14691] = 8'h57;
Memory[14690] = 8'h50;
Memory[14689] = 8'h40;
Memory[14688] = 8'h6F;
Memory[14695] = 8'h0E;
Memory[14694] = 8'h0C;
Memory[14693] = 8'hA2;
Memory[14692] = 8'h03;
Memory[14699] = 8'h00;
Memory[14698] = 8'h32;
Memory[14697] = 8'h22;
Memory[14696] = 8'hB3;
Memory[14703] = 8'h00;
Memory[14702] = 8'h02;
Memory[14701] = 8'h84;
Memory[14700] = 8'h63;
Memory[14707] = 8'h56;
Memory[14706] = 8'h90;
Memory[14705] = 8'h40;
Memory[14704] = 8'h6F;
Memory[14711] = 8'h0D;
Memory[14710] = 8'hCC;
Memory[14709] = 8'hA2;
Memory[14708] = 8'h03;
Memory[14715] = 8'h00;
Memory[14714] = 8'h32;
Memory[14713] = 8'h22;
Memory[14712] = 8'hB3;
Memory[14719] = 8'h00;
Memory[14718] = 8'h02;
Memory[14717] = 8'h84;
Memory[14716] = 8'h63;
Memory[14723] = 8'h55;
Memory[14722] = 8'hD0;
Memory[14721] = 8'h40;
Memory[14720] = 8'h6F;
Memory[14727] = 8'h0D;
Memory[14726] = 8'h8C;
Memory[14725] = 8'hA2;
Memory[14724] = 8'h03;
Memory[14731] = 8'h00;
Memory[14730] = 8'h32;
Memory[14729] = 8'h22;
Memory[14728] = 8'hB3;
Memory[14735] = 8'h00;
Memory[14734] = 8'h02;
Memory[14733] = 8'h84;
Memory[14732] = 8'h63;
Memory[14739] = 8'h55;
Memory[14738] = 8'h10;
Memory[14737] = 8'h40;
Memory[14736] = 8'h6F;
Memory[14743] = 8'h0D;
Memory[14742] = 8'h4C;
Memory[14741] = 8'hA2;
Memory[14740] = 8'h03;
Memory[14747] = 8'h00;
Memory[14746] = 8'h32;
Memory[14745] = 8'h22;
Memory[14744] = 8'hB3;
Memory[14751] = 8'h00;
Memory[14750] = 8'h02;
Memory[14749] = 8'h84;
Memory[14748] = 8'h63;
Memory[14755] = 8'h54;
Memory[14754] = 8'h50;
Memory[14753] = 8'h40;
Memory[14752] = 8'h6F;
Memory[14759] = 8'h0D;
Memory[14758] = 8'h0C;
Memory[14757] = 8'hA2;
Memory[14756] = 8'h03;
Memory[14763] = 8'h00;
Memory[14762] = 8'h32;
Memory[14761] = 8'h22;
Memory[14760] = 8'hB3;
Memory[14767] = 8'h00;
Memory[14766] = 8'h02;
Memory[14765] = 8'h84;
Memory[14764] = 8'h63;
Memory[14771] = 8'h53;
Memory[14770] = 8'h90;
Memory[14769] = 8'h40;
Memory[14768] = 8'h6F;
Memory[14775] = 8'h0C;
Memory[14774] = 8'hCC;
Memory[14773] = 8'hA2;
Memory[14772] = 8'h03;
Memory[14779] = 8'h00;
Memory[14778] = 8'h32;
Memory[14777] = 8'h22;
Memory[14776] = 8'hB3;
Memory[14783] = 8'h00;
Memory[14782] = 8'h02;
Memory[14781] = 8'h84;
Memory[14780] = 8'h63;
Memory[14787] = 8'h52;
Memory[14786] = 8'hD0;
Memory[14785] = 8'h40;
Memory[14784] = 8'h6F;
Memory[14791] = 8'h0C;
Memory[14790] = 8'h8C;
Memory[14789] = 8'hA2;
Memory[14788] = 8'h03;
Memory[14795] = 8'h00;
Memory[14794] = 8'h32;
Memory[14793] = 8'h22;
Memory[14792] = 8'hB3;
Memory[14799] = 8'h00;
Memory[14798] = 8'h02;
Memory[14797] = 8'h84;
Memory[14796] = 8'h63;
Memory[14803] = 8'h52;
Memory[14802] = 8'h10;
Memory[14801] = 8'h40;
Memory[14800] = 8'h6F;
Memory[14807] = 8'h0C;
Memory[14806] = 8'h4C;
Memory[14805] = 8'hA2;
Memory[14804] = 8'h03;
Memory[14811] = 8'h00;
Memory[14810] = 8'h32;
Memory[14809] = 8'h22;
Memory[14808] = 8'hB3;
Memory[14815] = 8'h00;
Memory[14814] = 8'h02;
Memory[14813] = 8'h84;
Memory[14812] = 8'h63;
Memory[14819] = 8'h51;
Memory[14818] = 8'h50;
Memory[14817] = 8'h40;
Memory[14816] = 8'h6F;
Memory[14823] = 8'h0C;
Memory[14822] = 8'h0C;
Memory[14821] = 8'hA2;
Memory[14820] = 8'h03;
Memory[14827] = 8'h00;
Memory[14826] = 8'h32;
Memory[14825] = 8'h22;
Memory[14824] = 8'hB3;
Memory[14831] = 8'h00;
Memory[14830] = 8'h02;
Memory[14829] = 8'h84;
Memory[14828] = 8'h63;
Memory[14835] = 8'h50;
Memory[14834] = 8'h90;
Memory[14833] = 8'h40;
Memory[14832] = 8'h6F;
Memory[14839] = 8'h0B;
Memory[14838] = 8'hCC;
Memory[14837] = 8'hA2;
Memory[14836] = 8'h03;
Memory[14843] = 8'h00;
Memory[14842] = 8'h32;
Memory[14841] = 8'h22;
Memory[14840] = 8'hB3;
Memory[14847] = 8'h00;
Memory[14846] = 8'h02;
Memory[14845] = 8'h84;
Memory[14844] = 8'h63;
Memory[14851] = 8'h4F;
Memory[14850] = 8'hD0;
Memory[14849] = 8'h40;
Memory[14848] = 8'h6F;
Memory[14855] = 8'h0B;
Memory[14854] = 8'h8C;
Memory[14853] = 8'hA2;
Memory[14852] = 8'h03;
Memory[14859] = 8'h00;
Memory[14858] = 8'h32;
Memory[14857] = 8'h22;
Memory[14856] = 8'hB3;
Memory[14863] = 8'h00;
Memory[14862] = 8'h02;
Memory[14861] = 8'h84;
Memory[14860] = 8'h63;
Memory[14867] = 8'h4F;
Memory[14866] = 8'h10;
Memory[14865] = 8'h40;
Memory[14864] = 8'h6F;
Memory[14871] = 8'h0B;
Memory[14870] = 8'h4C;
Memory[14869] = 8'hA2;
Memory[14868] = 8'h03;
Memory[14875] = 8'h00;
Memory[14874] = 8'h32;
Memory[14873] = 8'h22;
Memory[14872] = 8'hB3;
Memory[14879] = 8'h00;
Memory[14878] = 8'h02;
Memory[14877] = 8'h84;
Memory[14876] = 8'h63;
Memory[14883] = 8'h4E;
Memory[14882] = 8'h50;
Memory[14881] = 8'h40;
Memory[14880] = 8'h6F;
Memory[14887] = 8'h0B;
Memory[14886] = 8'h0C;
Memory[14885] = 8'hA2;
Memory[14884] = 8'h03;
Memory[14891] = 8'h00;
Memory[14890] = 8'h32;
Memory[14889] = 8'h22;
Memory[14888] = 8'hB3;
Memory[14895] = 8'h00;
Memory[14894] = 8'h02;
Memory[14893] = 8'h84;
Memory[14892] = 8'h63;
Memory[14899] = 8'h4D;
Memory[14898] = 8'h90;
Memory[14897] = 8'h40;
Memory[14896] = 8'h6F;
Memory[14903] = 8'h0A;
Memory[14902] = 8'hCC;
Memory[14901] = 8'hA2;
Memory[14900] = 8'h03;
Memory[14907] = 8'h00;
Memory[14906] = 8'h32;
Memory[14905] = 8'h22;
Memory[14904] = 8'hB3;
Memory[14911] = 8'h00;
Memory[14910] = 8'h02;
Memory[14909] = 8'h84;
Memory[14908] = 8'h63;
Memory[14915] = 8'h4C;
Memory[14914] = 8'hD0;
Memory[14913] = 8'h40;
Memory[14912] = 8'h6F;
Memory[14919] = 8'h0A;
Memory[14918] = 8'h8C;
Memory[14917] = 8'hA2;
Memory[14916] = 8'h03;
Memory[14923] = 8'h00;
Memory[14922] = 8'h32;
Memory[14921] = 8'h22;
Memory[14920] = 8'hB3;
Memory[14927] = 8'h00;
Memory[14926] = 8'h02;
Memory[14925] = 8'h84;
Memory[14924] = 8'h63;
Memory[14931] = 8'h4C;
Memory[14930] = 8'h10;
Memory[14929] = 8'h40;
Memory[14928] = 8'h6F;
Memory[14935] = 8'h0A;
Memory[14934] = 8'h4C;
Memory[14933] = 8'hA2;
Memory[14932] = 8'h03;
Memory[14939] = 8'h00;
Memory[14938] = 8'h32;
Memory[14937] = 8'h22;
Memory[14936] = 8'hB3;
Memory[14943] = 8'h00;
Memory[14942] = 8'h02;
Memory[14941] = 8'h84;
Memory[14940] = 8'h63;
Memory[14947] = 8'h4B;
Memory[14946] = 8'h50;
Memory[14945] = 8'h40;
Memory[14944] = 8'h6F;
Memory[14951] = 8'h0A;
Memory[14950] = 8'h0C;
Memory[14949] = 8'hA2;
Memory[14948] = 8'h03;
Memory[14955] = 8'h00;
Memory[14954] = 8'h32;
Memory[14953] = 8'h22;
Memory[14952] = 8'hB3;
Memory[14959] = 8'h00;
Memory[14958] = 8'h02;
Memory[14957] = 8'h84;
Memory[14956] = 8'h63;
Memory[14963] = 8'h4A;
Memory[14962] = 8'h90;
Memory[14961] = 8'h40;
Memory[14960] = 8'h6F;
Memory[14967] = 8'h09;
Memory[14966] = 8'hCC;
Memory[14965] = 8'hA2;
Memory[14964] = 8'h03;
Memory[14971] = 8'h00;
Memory[14970] = 8'h32;
Memory[14969] = 8'h22;
Memory[14968] = 8'hB3;
Memory[14975] = 8'h00;
Memory[14974] = 8'h02;
Memory[14973] = 8'h84;
Memory[14972] = 8'h63;
Memory[14979] = 8'h49;
Memory[14978] = 8'hD0;
Memory[14977] = 8'h40;
Memory[14976] = 8'h6F;
Memory[14983] = 8'h09;
Memory[14982] = 8'h8C;
Memory[14981] = 8'hA2;
Memory[14980] = 8'h03;
Memory[14987] = 8'h00;
Memory[14986] = 8'h32;
Memory[14985] = 8'h22;
Memory[14984] = 8'hB3;
Memory[14991] = 8'h00;
Memory[14990] = 8'h02;
Memory[14989] = 8'h84;
Memory[14988] = 8'h63;
Memory[14995] = 8'h49;
Memory[14994] = 8'h10;
Memory[14993] = 8'h40;
Memory[14992] = 8'h6F;
Memory[14999] = 8'h09;
Memory[14998] = 8'h4C;
Memory[14997] = 8'hA2;
Memory[14996] = 8'h03;
Memory[15003] = 8'h00;
Memory[15002] = 8'h32;
Memory[15001] = 8'h22;
Memory[15000] = 8'hB3;
Memory[15007] = 8'h00;
Memory[15006] = 8'h02;
Memory[15005] = 8'h84;
Memory[15004] = 8'h63;
Memory[15011] = 8'h48;
Memory[15010] = 8'h50;
Memory[15009] = 8'h40;
Memory[15008] = 8'h6F;
Memory[15015] = 8'h09;
Memory[15014] = 8'h0C;
Memory[15013] = 8'hA2;
Memory[15012] = 8'h03;
Memory[15019] = 8'h00;
Memory[15018] = 8'h32;
Memory[15017] = 8'h22;
Memory[15016] = 8'hB3;
Memory[15023] = 8'h00;
Memory[15022] = 8'h02;
Memory[15021] = 8'h84;
Memory[15020] = 8'h63;
Memory[15027] = 8'h47;
Memory[15026] = 8'h90;
Memory[15025] = 8'h40;
Memory[15024] = 8'h6F;
Memory[15031] = 8'h08;
Memory[15030] = 8'hCC;
Memory[15029] = 8'hA2;
Memory[15028] = 8'h03;
Memory[15035] = 8'h00;
Memory[15034] = 8'h32;
Memory[15033] = 8'h22;
Memory[15032] = 8'hB3;
Memory[15039] = 8'h00;
Memory[15038] = 8'h02;
Memory[15037] = 8'h84;
Memory[15036] = 8'h63;
Memory[15043] = 8'h46;
Memory[15042] = 8'hD0;
Memory[15041] = 8'h40;
Memory[15040] = 8'h6F;
Memory[15047] = 8'h08;
Memory[15046] = 8'h8C;
Memory[15045] = 8'hA2;
Memory[15044] = 8'h03;
Memory[15051] = 8'h00;
Memory[15050] = 8'h32;
Memory[15049] = 8'h22;
Memory[15048] = 8'hB3;
Memory[15055] = 8'h00;
Memory[15054] = 8'h02;
Memory[15053] = 8'h84;
Memory[15052] = 8'h63;
Memory[15059] = 8'h46;
Memory[15058] = 8'h10;
Memory[15057] = 8'h40;
Memory[15056] = 8'h6F;
Memory[15063] = 8'h08;
Memory[15062] = 8'h4C;
Memory[15061] = 8'hA2;
Memory[15060] = 8'h03;
Memory[15067] = 8'h00;
Memory[15066] = 8'h32;
Memory[15065] = 8'h22;
Memory[15064] = 8'hB3;
Memory[15071] = 8'h00;
Memory[15070] = 8'h02;
Memory[15069] = 8'h84;
Memory[15068] = 8'h63;
Memory[15075] = 8'h45;
Memory[15074] = 8'h50;
Memory[15073] = 8'h40;
Memory[15072] = 8'h6F;
Memory[15079] = 8'h08;
Memory[15078] = 8'h0C;
Memory[15077] = 8'hA2;
Memory[15076] = 8'h03;
Memory[15083] = 8'h00;
Memory[15082] = 8'h32;
Memory[15081] = 8'h22;
Memory[15080] = 8'hB3;
Memory[15087] = 8'h00;
Memory[15086] = 8'h02;
Memory[15085] = 8'h84;
Memory[15084] = 8'h63;
Memory[15091] = 8'h44;
Memory[15090] = 8'h90;
Memory[15089] = 8'h40;
Memory[15088] = 8'h6F;
Memory[15095] = 8'h07;
Memory[15094] = 8'hCC;
Memory[15093] = 8'hA2;
Memory[15092] = 8'h03;
Memory[15099] = 8'h00;
Memory[15098] = 8'h32;
Memory[15097] = 8'h22;
Memory[15096] = 8'hB3;
Memory[15103] = 8'h00;
Memory[15102] = 8'h02;
Memory[15101] = 8'h84;
Memory[15100] = 8'h63;
Memory[15107] = 8'h43;
Memory[15106] = 8'hD0;
Memory[15105] = 8'h40;
Memory[15104] = 8'h6F;
Memory[15111] = 8'h07;
Memory[15110] = 8'h8C;
Memory[15109] = 8'hA2;
Memory[15108] = 8'h03;
Memory[15115] = 8'h00;
Memory[15114] = 8'h32;
Memory[15113] = 8'h22;
Memory[15112] = 8'hB3;
Memory[15119] = 8'h00;
Memory[15118] = 8'h02;
Memory[15117] = 8'h84;
Memory[15116] = 8'h63;
Memory[15123] = 8'h43;
Memory[15122] = 8'h10;
Memory[15121] = 8'h40;
Memory[15120] = 8'h6F;
Memory[15127] = 8'h07;
Memory[15126] = 8'h4C;
Memory[15125] = 8'hA2;
Memory[15124] = 8'h03;
Memory[15131] = 8'h00;
Memory[15130] = 8'h32;
Memory[15129] = 8'h22;
Memory[15128] = 8'hB3;
Memory[15135] = 8'h00;
Memory[15134] = 8'h02;
Memory[15133] = 8'h84;
Memory[15132] = 8'h63;
Memory[15139] = 8'h42;
Memory[15138] = 8'h50;
Memory[15137] = 8'h40;
Memory[15136] = 8'h6F;
Memory[15143] = 8'h07;
Memory[15142] = 8'h0C;
Memory[15141] = 8'hA2;
Memory[15140] = 8'h03;
Memory[15147] = 8'h00;
Memory[15146] = 8'h32;
Memory[15145] = 8'h22;
Memory[15144] = 8'hB3;
Memory[15151] = 8'h00;
Memory[15150] = 8'h02;
Memory[15149] = 8'h84;
Memory[15148] = 8'h63;
Memory[15155] = 8'h41;
Memory[15154] = 8'h90;
Memory[15153] = 8'h40;
Memory[15152] = 8'h6F;
Memory[15159] = 8'h06;
Memory[15158] = 8'hCC;
Memory[15157] = 8'hA2;
Memory[15156] = 8'h03;
Memory[15163] = 8'h00;
Memory[15162] = 8'h32;
Memory[15161] = 8'h22;
Memory[15160] = 8'hB3;
Memory[15167] = 8'h00;
Memory[15166] = 8'h02;
Memory[15165] = 8'h84;
Memory[15164] = 8'h63;
Memory[15171] = 8'h40;
Memory[15170] = 8'hD0;
Memory[15169] = 8'h40;
Memory[15168] = 8'h6F;
Memory[15175] = 8'h06;
Memory[15174] = 8'h8C;
Memory[15173] = 8'hA2;
Memory[15172] = 8'h03;
Memory[15179] = 8'h00;
Memory[15178] = 8'h32;
Memory[15177] = 8'h22;
Memory[15176] = 8'hB3;
Memory[15183] = 8'h00;
Memory[15182] = 8'h02;
Memory[15181] = 8'h84;
Memory[15180] = 8'h63;
Memory[15187] = 8'h40;
Memory[15186] = 8'h10;
Memory[15185] = 8'h40;
Memory[15184] = 8'h6F;
Memory[15191] = 8'h06;
Memory[15190] = 8'h4C;
Memory[15189] = 8'hA2;
Memory[15188] = 8'h03;
Memory[15195] = 8'h00;
Memory[15194] = 8'h32;
Memory[15193] = 8'h22;
Memory[15192] = 8'hB3;
Memory[15199] = 8'h00;
Memory[15198] = 8'h02;
Memory[15197] = 8'h84;
Memory[15196] = 8'h63;
Memory[15203] = 8'h3F;
Memory[15202] = 8'h50;
Memory[15201] = 8'h40;
Memory[15200] = 8'h6F;
Memory[15207] = 8'h06;
Memory[15206] = 8'h0C;
Memory[15205] = 8'hA2;
Memory[15204] = 8'h03;
Memory[15211] = 8'h00;
Memory[15210] = 8'h32;
Memory[15209] = 8'h22;
Memory[15208] = 8'hB3;
Memory[15215] = 8'h00;
Memory[15214] = 8'h02;
Memory[15213] = 8'h84;
Memory[15212] = 8'h63;
Memory[15219] = 8'h3E;
Memory[15218] = 8'h90;
Memory[15217] = 8'h40;
Memory[15216] = 8'h6F;
Memory[15223] = 8'h05;
Memory[15222] = 8'hCC;
Memory[15221] = 8'hA2;
Memory[15220] = 8'h03;
Memory[15227] = 8'h00;
Memory[15226] = 8'h32;
Memory[15225] = 8'h22;
Memory[15224] = 8'hB3;
Memory[15231] = 8'h00;
Memory[15230] = 8'h02;
Memory[15229] = 8'h84;
Memory[15228] = 8'h63;
Memory[15235] = 8'h3D;
Memory[15234] = 8'hD0;
Memory[15233] = 8'h40;
Memory[15232] = 8'h6F;
Memory[15239] = 8'h05;
Memory[15238] = 8'h8C;
Memory[15237] = 8'hA2;
Memory[15236] = 8'h03;
Memory[15243] = 8'h00;
Memory[15242] = 8'h32;
Memory[15241] = 8'h22;
Memory[15240] = 8'hB3;
Memory[15247] = 8'h00;
Memory[15246] = 8'h02;
Memory[15245] = 8'h84;
Memory[15244] = 8'h63;
Memory[15251] = 8'h3D;
Memory[15250] = 8'h10;
Memory[15249] = 8'h40;
Memory[15248] = 8'h6F;
Memory[15255] = 8'h05;
Memory[15254] = 8'h4C;
Memory[15253] = 8'hA2;
Memory[15252] = 8'h03;
Memory[15259] = 8'h00;
Memory[15258] = 8'h32;
Memory[15257] = 8'h22;
Memory[15256] = 8'hB3;
Memory[15263] = 8'h00;
Memory[15262] = 8'h02;
Memory[15261] = 8'h84;
Memory[15260] = 8'h63;
Memory[15267] = 8'h3C;
Memory[15266] = 8'h50;
Memory[15265] = 8'h40;
Memory[15264] = 8'h6F;
Memory[15271] = 8'h05;
Memory[15270] = 8'h0C;
Memory[15269] = 8'hA2;
Memory[15268] = 8'h03;
Memory[15275] = 8'h00;
Memory[15274] = 8'h32;
Memory[15273] = 8'h22;
Memory[15272] = 8'hB3;
Memory[15279] = 8'h00;
Memory[15278] = 8'h02;
Memory[15277] = 8'h84;
Memory[15276] = 8'h63;
Memory[15283] = 8'h3B;
Memory[15282] = 8'h90;
Memory[15281] = 8'h40;
Memory[15280] = 8'h6F;
Memory[15287] = 8'h04;
Memory[15286] = 8'hCC;
Memory[15285] = 8'hA2;
Memory[15284] = 8'h03;
Memory[15291] = 8'h00;
Memory[15290] = 8'h32;
Memory[15289] = 8'h22;
Memory[15288] = 8'hB3;
Memory[15295] = 8'h00;
Memory[15294] = 8'h02;
Memory[15293] = 8'h84;
Memory[15292] = 8'h63;
Memory[15299] = 8'h3A;
Memory[15298] = 8'hD0;
Memory[15297] = 8'h40;
Memory[15296] = 8'h6F;
Memory[15303] = 8'h04;
Memory[15302] = 8'h8C;
Memory[15301] = 8'hA2;
Memory[15300] = 8'h03;
Memory[15307] = 8'h00;
Memory[15306] = 8'h32;
Memory[15305] = 8'h22;
Memory[15304] = 8'hB3;
Memory[15311] = 8'h00;
Memory[15310] = 8'h02;
Memory[15309] = 8'h84;
Memory[15308] = 8'h63;
Memory[15315] = 8'h3A;
Memory[15314] = 8'h10;
Memory[15313] = 8'h40;
Memory[15312] = 8'h6F;
Memory[15319] = 8'h04;
Memory[15318] = 8'h4C;
Memory[15317] = 8'hA2;
Memory[15316] = 8'h03;
Memory[15323] = 8'h00;
Memory[15322] = 8'h32;
Memory[15321] = 8'h22;
Memory[15320] = 8'hB3;
Memory[15327] = 8'h00;
Memory[15326] = 8'h02;
Memory[15325] = 8'h84;
Memory[15324] = 8'h63;
Memory[15331] = 8'h39;
Memory[15330] = 8'h50;
Memory[15329] = 8'h40;
Memory[15328] = 8'h6F;
Memory[15335] = 8'h04;
Memory[15334] = 8'h0C;
Memory[15333] = 8'hA2;
Memory[15332] = 8'h03;
Memory[15339] = 8'h00;
Memory[15338] = 8'h32;
Memory[15337] = 8'h22;
Memory[15336] = 8'hB3;
Memory[15343] = 8'h00;
Memory[15342] = 8'h02;
Memory[15341] = 8'h84;
Memory[15340] = 8'h63;
Memory[15347] = 8'h38;
Memory[15346] = 8'h90;
Memory[15345] = 8'h40;
Memory[15344] = 8'h6F;
Memory[15351] = 8'h03;
Memory[15350] = 8'hCC;
Memory[15349] = 8'hA2;
Memory[15348] = 8'h03;
Memory[15355] = 8'h00;
Memory[15354] = 8'h32;
Memory[15353] = 8'h22;
Memory[15352] = 8'hB3;
Memory[15359] = 8'h00;
Memory[15358] = 8'h02;
Memory[15357] = 8'h84;
Memory[15356] = 8'h63;
Memory[15363] = 8'h37;
Memory[15362] = 8'hD0;
Memory[15361] = 8'h40;
Memory[15360] = 8'h6F;
Memory[15367] = 8'h03;
Memory[15366] = 8'h8C;
Memory[15365] = 8'hA2;
Memory[15364] = 8'h03;
Memory[15371] = 8'h00;
Memory[15370] = 8'h32;
Memory[15369] = 8'h22;
Memory[15368] = 8'hB3;
Memory[15375] = 8'h00;
Memory[15374] = 8'h02;
Memory[15373] = 8'h84;
Memory[15372] = 8'h63;
Memory[15379] = 8'h37;
Memory[15378] = 8'h10;
Memory[15377] = 8'h40;
Memory[15376] = 8'h6F;
Memory[15383] = 8'h03;
Memory[15382] = 8'h4C;
Memory[15381] = 8'hA2;
Memory[15380] = 8'h03;
Memory[15387] = 8'h00;
Memory[15386] = 8'h32;
Memory[15385] = 8'h22;
Memory[15384] = 8'hB3;
Memory[15391] = 8'h00;
Memory[15390] = 8'h02;
Memory[15389] = 8'h84;
Memory[15388] = 8'h63;
Memory[15395] = 8'h36;
Memory[15394] = 8'h50;
Memory[15393] = 8'h40;
Memory[15392] = 8'h6F;
Memory[15399] = 8'h03;
Memory[15398] = 8'h0C;
Memory[15397] = 8'hA2;
Memory[15396] = 8'h03;
Memory[15403] = 8'h00;
Memory[15402] = 8'h32;
Memory[15401] = 8'h22;
Memory[15400] = 8'hB3;
Memory[15407] = 8'h00;
Memory[15406] = 8'h02;
Memory[15405] = 8'h84;
Memory[15404] = 8'h63;
Memory[15411] = 8'h35;
Memory[15410] = 8'h90;
Memory[15409] = 8'h40;
Memory[15408] = 8'h6F;
Memory[15415] = 8'h02;
Memory[15414] = 8'hCC;
Memory[15413] = 8'hA2;
Memory[15412] = 8'h03;
Memory[15419] = 8'h00;
Memory[15418] = 8'h32;
Memory[15417] = 8'h22;
Memory[15416] = 8'hB3;
Memory[15423] = 8'h00;
Memory[15422] = 8'h02;
Memory[15421] = 8'h84;
Memory[15420] = 8'h63;
Memory[15427] = 8'h34;
Memory[15426] = 8'hD0;
Memory[15425] = 8'h40;
Memory[15424] = 8'h6F;
Memory[15431] = 8'h02;
Memory[15430] = 8'h8C;
Memory[15429] = 8'hA2;
Memory[15428] = 8'h03;
Memory[15435] = 8'h00;
Memory[15434] = 8'h32;
Memory[15433] = 8'h22;
Memory[15432] = 8'hB3;
Memory[15439] = 8'h00;
Memory[15438] = 8'h02;
Memory[15437] = 8'h84;
Memory[15436] = 8'h63;
Memory[15443] = 8'h34;
Memory[15442] = 8'h10;
Memory[15441] = 8'h40;
Memory[15440] = 8'h6F;
Memory[15447] = 8'h02;
Memory[15446] = 8'h4C;
Memory[15445] = 8'hA2;
Memory[15444] = 8'h03;
Memory[15451] = 8'h00;
Memory[15450] = 8'h32;
Memory[15449] = 8'h22;
Memory[15448] = 8'hB3;
Memory[15455] = 8'h00;
Memory[15454] = 8'h02;
Memory[15453] = 8'h84;
Memory[15452] = 8'h63;
Memory[15459] = 8'h33;
Memory[15458] = 8'h50;
Memory[15457] = 8'h40;
Memory[15456] = 8'h6F;
Memory[15463] = 8'h02;
Memory[15462] = 8'h0C;
Memory[15461] = 8'hA2;
Memory[15460] = 8'h03;
Memory[15467] = 8'h00;
Memory[15466] = 8'h32;
Memory[15465] = 8'h22;
Memory[15464] = 8'hB3;
Memory[15471] = 8'h00;
Memory[15470] = 8'h02;
Memory[15469] = 8'h84;
Memory[15468] = 8'h63;
Memory[15475] = 8'h32;
Memory[15474] = 8'h90;
Memory[15473] = 8'h40;
Memory[15472] = 8'h6F;
Memory[15479] = 8'h01;
Memory[15478] = 8'hCC;
Memory[15477] = 8'hA2;
Memory[15476] = 8'h03;
Memory[15483] = 8'h00;
Memory[15482] = 8'h32;
Memory[15481] = 8'h22;
Memory[15480] = 8'hB3;
Memory[15487] = 8'h00;
Memory[15486] = 8'h02;
Memory[15485] = 8'h84;
Memory[15484] = 8'h63;
Memory[15491] = 8'h31;
Memory[15490] = 8'hD0;
Memory[15489] = 8'h40;
Memory[15488] = 8'h6F;
Memory[15495] = 8'h01;
Memory[15494] = 8'h8C;
Memory[15493] = 8'hA2;
Memory[15492] = 8'h03;
Memory[15499] = 8'h00;
Memory[15498] = 8'h32;
Memory[15497] = 8'h22;
Memory[15496] = 8'hB3;
Memory[15503] = 8'h00;
Memory[15502] = 8'h02;
Memory[15501] = 8'h84;
Memory[15500] = 8'h63;
Memory[15507] = 8'h31;
Memory[15506] = 8'h10;
Memory[15505] = 8'h40;
Memory[15504] = 8'h6F;
Memory[15511] = 8'h01;
Memory[15510] = 8'h4C;
Memory[15509] = 8'hA2;
Memory[15508] = 8'h03;
Memory[15515] = 8'h00;
Memory[15514] = 8'h32;
Memory[15513] = 8'h22;
Memory[15512] = 8'hB3;
Memory[15519] = 8'h00;
Memory[15518] = 8'h02;
Memory[15517] = 8'h84;
Memory[15516] = 8'h63;
Memory[15523] = 8'h30;
Memory[15522] = 8'h50;
Memory[15521] = 8'h40;
Memory[15520] = 8'h6F;
Memory[15527] = 8'h01;
Memory[15526] = 8'h0C;
Memory[15525] = 8'hA2;
Memory[15524] = 8'h03;
Memory[15531] = 8'h00;
Memory[15530] = 8'h32;
Memory[15529] = 8'h22;
Memory[15528] = 8'hB3;
Memory[15535] = 8'h00;
Memory[15534] = 8'h02;
Memory[15533] = 8'h84;
Memory[15532] = 8'h63;
Memory[15539] = 8'h2F;
Memory[15538] = 8'h90;
Memory[15537] = 8'h40;
Memory[15536] = 8'h6F;
Memory[15543] = 8'h00;
Memory[15542] = 8'hCC;
Memory[15541] = 8'hA2;
Memory[15540] = 8'h03;
Memory[15547] = 8'h00;
Memory[15546] = 8'h32;
Memory[15545] = 8'h22;
Memory[15544] = 8'hB3;
Memory[15551] = 8'h00;
Memory[15550] = 8'h02;
Memory[15549] = 8'h84;
Memory[15548] = 8'h63;
Memory[15555] = 8'h2E;
Memory[15554] = 8'hD0;
Memory[15553] = 8'h40;
Memory[15552] = 8'h6F;
Memory[15559] = 8'h00;
Memory[15558] = 8'h8C;
Memory[15557] = 8'hA2;
Memory[15556] = 8'h03;
Memory[15563] = 8'h00;
Memory[15562] = 8'h32;
Memory[15561] = 8'h22;
Memory[15560] = 8'hB3;
Memory[15567] = 8'h00;
Memory[15566] = 8'h02;
Memory[15565] = 8'h84;
Memory[15564] = 8'h63;
Memory[15571] = 8'h2E;
Memory[15570] = 8'h10;
Memory[15569] = 8'h40;
Memory[15568] = 8'h6F;
Memory[15575] = 8'h00;
Memory[15574] = 8'h4C;
Memory[15573] = 8'hA2;
Memory[15572] = 8'h03;
Memory[15579] = 8'h00;
Memory[15578] = 8'h32;
Memory[15577] = 8'h22;
Memory[15576] = 8'hB3;
Memory[15583] = 8'h00;
Memory[15582] = 8'h02;
Memory[15581] = 8'h84;
Memory[15580] = 8'h63;
Memory[15587] = 8'h2D;
Memory[15586] = 8'h50;
Memory[15585] = 8'h40;
Memory[15584] = 8'h6F;
Memory[15591] = 8'h00;
Memory[15590] = 8'h0C;
Memory[15589] = 8'hA2;
Memory[15588] = 8'h03;
Memory[15595] = 8'h00;
Memory[15594] = 8'h32;
Memory[15593] = 8'h22;
Memory[15592] = 8'hB3;
Memory[15599] = 8'h00;
Memory[15598] = 8'h02;
Memory[15597] = 8'h84;
Memory[15596] = 8'h63;
Memory[15603] = 8'h2C;
Memory[15602] = 8'h90;
Memory[15601] = 8'h40;
Memory[15600] = 8'h6F;
Memory[15607] = 8'h12;
Memory[15606] = 8'h40;
Memory[15605] = 8'h20;
Memory[15604] = 8'h6F;
Memory[15611] = 8'h00;
Memory[15610] = 8'h00;
Memory[15609] = 8'h00;
Memory[15608] = 8'h00;
Memory[15615] = 8'h00;
Memory[15614] = 8'h00;
Memory[15613] = 8'h03;
Memory[15612] = 8'hE8;
Memory[15619] = 8'h00;
Memory[15618] = 8'h00;
Memory[15617] = 8'h07;
Memory[15616] = 8'hD0;
Memory[15623] = 8'h00;
Memory[15622] = 8'h00;
Memory[15621] = 8'h0B;
Memory[15620] = 8'hB8;
Memory[15627] = 8'h00;
Memory[15626] = 8'h00;
Memory[15625] = 8'h0F;
Memory[15624] = 8'hA0;
Memory[15631] = 8'h00;
Memory[15630] = 8'h00;
Memory[15629] = 8'h13;
Memory[15628] = 8'h88;
Memory[15635] = 8'h00;
Memory[15634] = 8'h00;
Memory[15633] = 8'h17;
Memory[15632] = 8'h70;
Memory[15639] = 8'h00;
Memory[15638] = 8'h00;
Memory[15637] = 8'h1B;
Memory[15636] = 8'h58;
Memory[15643] = 8'h00;
Memory[15642] = 8'h00;
Memory[15641] = 8'h1F;
Memory[15640] = 8'h40;
Memory[15647] = 8'h00;
Memory[15646] = 8'h00;
Memory[15645] = 8'h23;
Memory[15644] = 8'h28;
Memory[15651] = 8'h00;
Memory[15650] = 8'h00;
Memory[15649] = 8'h27;
Memory[15648] = 8'h10;
Memory[15655] = 8'h00;
Memory[15654] = 8'h00;
Memory[15653] = 8'h2A;
Memory[15652] = 8'hF8;
Memory[15659] = 8'h00;
Memory[15658] = 8'h00;
Memory[15657] = 8'h2E;
Memory[15656] = 8'hE0;
Memory[15663] = 8'h00;
Memory[15662] = 8'h00;
Memory[15661] = 8'h32;
Memory[15660] = 8'hC8;
Memory[15667] = 8'h00;
Memory[15666] = 8'h00;
Memory[15665] = 8'h36;
Memory[15664] = 8'hB0;
Memory[15671] = 8'h00;
Memory[15670] = 8'h00;
Memory[15669] = 8'h3A;
Memory[15668] = 8'h98;
Memory[15675] = 8'h00;
Memory[15674] = 8'h00;
Memory[15673] = 8'h3E;
Memory[15672] = 8'h80;
Memory[15679] = 8'h00;
Memory[15678] = 8'h00;
Memory[15677] = 8'h42;
Memory[15676] = 8'h68;
Memory[15683] = 8'h00;
Memory[15682] = 8'h00;
Memory[15681] = 8'h46;
Memory[15680] = 8'h50;
Memory[15687] = 8'h00;
Memory[15686] = 8'h00;
Memory[15685] = 8'h4A;
Memory[15684] = 8'h38;
Memory[15691] = 8'h00;
Memory[15690] = 8'h00;
Memory[15689] = 8'h4E;
Memory[15688] = 8'h20;
Memory[15695] = 8'h00;
Memory[15694] = 8'h00;
Memory[15693] = 8'h52;
Memory[15692] = 8'h08;
Memory[15699] = 8'h00;
Memory[15698] = 8'h00;
Memory[15697] = 8'h55;
Memory[15696] = 8'hF0;
Memory[15703] = 8'h00;
Memory[15702] = 8'h00;
Memory[15701] = 8'h59;
Memory[15700] = 8'hD8;
Memory[15707] = 8'h00;
Memory[15706] = 8'h00;
Memory[15705] = 8'h5D;
Memory[15704] = 8'hC0;
Memory[15711] = 8'h00;
Memory[15710] = 8'h00;
Memory[15709] = 8'h5F;
Memory[15708] = 8'hB4;
Memory[15715] = 8'h00;
Memory[15714] = 8'h00;
Memory[15713] = 8'h61;
Memory[15712] = 8'hA8;
Memory[15719] = 8'h00;
Memory[15718] = 8'h00;
Memory[15717] = 8'h63;
Memory[15716] = 8'h9C;
Memory[15723] = 8'h00;
Memory[15722] = 8'h00;
Memory[15721] = 8'h65;
Memory[15720] = 8'h90;
Memory[15727] = 8'h00;
Memory[15726] = 8'h00;
Memory[15725] = 8'h67;
Memory[15724] = 8'h84;
Memory[15731] = 8'h00;
Memory[15730] = 8'h00;
Memory[15729] = 8'h69;
Memory[15728] = 8'h78;
Memory[15735] = 8'h00;
Memory[15734] = 8'h00;
Memory[15733] = 8'h6B;
Memory[15732] = 8'h6C;
Memory[15739] = 8'h00;
Memory[15738] = 8'h00;
Memory[15737] = 8'h6D;
Memory[15736] = 8'h60;
Memory[15743] = 8'h00;
Memory[15742] = 8'h00;
Memory[15741] = 8'h6F;
Memory[15740] = 8'h54;
Memory[15747] = 8'h00;
Memory[15746] = 8'h00;
Memory[15745] = 8'h71;
Memory[15744] = 8'h48;
Memory[15751] = 8'h00;
Memory[15750] = 8'h00;
Memory[15749] = 8'h73;
Memory[15748] = 8'h3C;
Memory[15755] = 8'h00;
Memory[15754] = 8'h00;
Memory[15753] = 8'h75;
Memory[15752] = 8'h30;
Memory[15759] = 8'h00;
Memory[15758] = 8'h00;
Memory[15757] = 8'h77;
Memory[15756] = 8'h24;
Memory[15763] = 8'h00;
Memory[15762] = 8'h00;
Memory[15761] = 8'h79;
Memory[15760] = 8'h18;
Memory[15767] = 8'h00;
Memory[15766] = 8'h00;
Memory[15765] = 8'h7B;
Memory[15764] = 8'h0C;
Memory[15771] = 8'h00;
Memory[15770] = 8'h00;
Memory[15769] = 8'h7D;
Memory[15768] = 8'h00;
Memory[15775] = 8'h00;
Memory[15774] = 8'h00;
Memory[15773] = 8'h7E;
Memory[15772] = 8'hF4;
Memory[15779] = 8'h00;
Memory[15778] = 8'h00;
Memory[15777] = 8'h80;
Memory[15776] = 8'hE8;
Memory[15783] = 8'h00;
Memory[15782] = 8'h00;
Memory[15781] = 8'h82;
Memory[15780] = 8'hDC;
Memory[15787] = 8'h00;
Memory[15786] = 8'h00;
Memory[15785] = 8'h84;
Memory[15784] = 8'hD0;
Memory[15791] = 8'h00;
Memory[15790] = 8'h00;
Memory[15789] = 8'h86;
Memory[15788] = 8'hC4;
Memory[15795] = 8'h00;
Memory[15794] = 8'h00;
Memory[15793] = 8'h88;
Memory[15792] = 8'hB8;
Memory[15799] = 8'h00;
Memory[15798] = 8'h00;
Memory[15797] = 8'h8A;
Memory[15796] = 8'hAC;
Memory[15803] = 8'h00;
Memory[15802] = 8'h00;
Memory[15801] = 8'h8C;
Memory[15800] = 8'hA0;
Memory[15807] = 8'h00;
Memory[15806] = 8'h00;
Memory[15805] = 8'h8E;
Memory[15804] = 8'h94;
Memory[15811] = 8'h00;
Memory[15810] = 8'h00;
Memory[15809] = 8'h90;
Memory[15808] = 8'h88;
Memory[15815] = 8'h00;
Memory[15814] = 8'h00;
Memory[15813] = 8'h92;
Memory[15812] = 8'h7C;
Memory[15819] = 8'h00;
Memory[15818] = 8'h00;
Memory[15817] = 8'h94;
Memory[15816] = 8'h70;
Memory[15823] = 8'h00;
Memory[15822] = 8'h00;
Memory[15821] = 8'h96;
Memory[15820] = 8'h64;
Memory[15827] = 8'h00;
Memory[15826] = 8'h00;
Memory[15825] = 8'h9B;
Memory[15824] = 8'h46;
Memory[15831] = 8'h00;
Memory[15830] = 8'h00;
Memory[15829] = 8'h9C;
Memory[15828] = 8'h40;
Memory[15835] = 8'h00;
Memory[15834] = 8'h00;
Memory[15833] = 8'h9D;
Memory[15832] = 8'h3A;
Memory[15839] = 8'h00;
Memory[15838] = 8'h00;
Memory[15837] = 8'h9E;
Memory[15836] = 8'h34;
Memory[15843] = 8'h00;
Memory[15842] = 8'h00;
Memory[15841] = 8'h9F;
Memory[15840] = 8'h2E;
Memory[15847] = 8'h00;
Memory[15846] = 8'h00;
Memory[15845] = 8'hA0;
Memory[15844] = 8'h28;
Memory[15851] = 8'h00;
Memory[15850] = 8'h00;
Memory[15849] = 8'hA1;
Memory[15848] = 8'h22;
Memory[15855] = 8'h00;
Memory[15854] = 8'h00;
Memory[15853] = 8'hA2;
Memory[15852] = 8'h1C;
Memory[15859] = 8'h00;
Memory[15858] = 8'h00;
Memory[15857] = 8'hA3;
Memory[15856] = 8'h16;
Memory[15863] = 8'h00;
Memory[15862] = 8'h00;
Memory[15861] = 8'hA4;
Memory[15860] = 8'h10;
Memory[15867] = 8'h00;
Memory[15866] = 8'h00;
Memory[15865] = 8'hA5;
Memory[15864] = 8'h0A;
Memory[15871] = 8'h00;
Memory[15870] = 8'h00;
Memory[15869] = 8'hA6;
Memory[15868] = 8'h04;
Memory[15875] = 8'h00;
Memory[15874] = 8'h00;
Memory[15873] = 8'hA6;
Memory[15872] = 8'hFE;
Memory[15879] = 8'h00;
Memory[15878] = 8'h00;
Memory[15877] = 8'hA7;
Memory[15876] = 8'hF8;
Memory[15883] = 8'h00;
Memory[15882] = 8'h00;
Memory[15881] = 8'hA8;
Memory[15880] = 8'hF2;
Memory[15887] = 8'h00;
Memory[15886] = 8'h00;
Memory[15885] = 8'hA9;
Memory[15884] = 8'hEC;
Memory[15891] = 8'h00;
Memory[15890] = 8'h00;
Memory[15889] = 8'hAA;
Memory[15888] = 8'hE6;
Memory[15895] = 8'h00;
Memory[15894] = 8'h00;
Memory[15893] = 8'hAB;
Memory[15892] = 8'hE0;
Memory[15899] = 8'h00;
Memory[15898] = 8'h00;
Memory[15897] = 8'hAC;
Memory[15896] = 8'hDA;
Memory[15903] = 8'h00;
Memory[15902] = 8'h00;
Memory[15901] = 8'hAD;
Memory[15900] = 8'hD4;
Memory[15907] = 8'h00;
Memory[15906] = 8'h00;
Memory[15905] = 8'hAE;
Memory[15904] = 8'hCE;
Memory[15911] = 8'h00;
Memory[15910] = 8'h00;
Memory[15909] = 8'hAF;
Memory[15908] = 8'hC8;
Memory[15915] = 8'h00;
Memory[15914] = 8'h00;
Memory[15913] = 8'hB0;
Memory[15912] = 8'hC2;
Memory[15919] = 8'h00;
Memory[15918] = 8'h00;
Memory[15917] = 8'hB1;
Memory[15916] = 8'hBC;
Memory[15923] = 8'h00;
Memory[15922] = 8'h00;
Memory[15921] = 8'hB2;
Memory[15920] = 8'hB6;
Memory[15927] = 8'h00;
Memory[15926] = 8'h00;
Memory[15925] = 8'hB3;
Memory[15924] = 8'hB0;
Memory[15931] = 8'h00;
Memory[15930] = 8'h00;
Memory[15929] = 8'hB4;
Memory[15928] = 8'hAA;
Memory[15935] = 8'h00;
Memory[15934] = 8'h00;
Memory[15933] = 8'hB5;
Memory[15932] = 8'hA4;
Memory[15939] = 8'h00;
Memory[15938] = 8'h00;
Memory[15937] = 8'hB6;
Memory[15936] = 8'h9E;
Memory[15943] = 8'h00;
Memory[15942] = 8'h00;
Memory[15941] = 8'hB7;
Memory[15940] = 8'h98;
Memory[15947] = 8'h00;
Memory[15946] = 8'h00;
Memory[15945] = 8'hB8;
Memory[15944] = 8'h92;
Memory[15951] = 8'h00;
Memory[15950] = 8'h00;
Memory[15949] = 8'hB9;
Memory[15948] = 8'h8C;
Memory[15955] = 8'h00;
Memory[15954] = 8'h00;
Memory[15953] = 8'hBA;
Memory[15952] = 8'h86;
Memory[15959] = 8'h00;
Memory[15958] = 8'h00;
Memory[15957] = 8'hBB;
Memory[15956] = 8'h80;
Memory[15963] = 8'h00;
Memory[15962] = 8'h00;
Memory[15961] = 8'hBC;
Memory[15960] = 8'h7A;
Memory[15967] = 8'h00;
Memory[15966] = 8'h00;
Memory[15965] = 8'hBD;
Memory[15964] = 8'h74;
Memory[15971] = 8'h00;
Memory[15970] = 8'h00;
Memory[15969] = 8'hBE;
Memory[15968] = 8'h6E;
Memory[15975] = 8'h00;
Memory[15974] = 8'h00;
Memory[15973] = 8'hBF;
Memory[15972] = 8'h68;
Memory[15979] = 8'h00;
Memory[15978] = 8'h00;
Memory[15977] = 8'hC0;
Memory[15976] = 8'h62;
Memory[15983] = 8'h00;
Memory[15982] = 8'h00;
Memory[15981] = 8'hC1;
Memory[15980] = 8'h5C;
Memory[15987] = 8'h00;
Memory[15986] = 8'h00;
Memory[15985] = 8'hC2;
Memory[15984] = 8'h56;
Memory[15991] = 8'h00;
Memory[15990] = 8'h00;
Memory[15989] = 8'hC3;
Memory[15988] = 8'h50;
Memory[15995] = 8'h00;
Memory[15994] = 8'h00;
Memory[15993] = 8'hC4;
Memory[15992] = 8'h4A;
Memory[15999] = 8'h00;
Memory[15998] = 8'h00;
Memory[15997] = 8'hC5;
Memory[15996] = 8'h44;
Memory[16003] = 8'h00;
Memory[16002] = 8'h00;
Memory[16001] = 8'hC6;
Memory[16000] = 8'h3E;
Memory[16007] = 8'h00;
Memory[16006] = 8'h00;
Memory[16005] = 8'hC7;
Memory[16004] = 8'h38;
Memory[16011] = 8'h00;
Memory[16010] = 8'h00;
Memory[16009] = 8'hC8;
Memory[16008] = 8'h32;
Memory[16015] = 8'h00;
Memory[16014] = 8'h00;
Memory[16013] = 8'hC9;
Memory[16012] = 8'h2C;
Memory[16019] = 8'h00;
Memory[16018] = 8'h00;
Memory[16017] = 8'hCA;
Memory[16016] = 8'h26;
Memory[16023] = 8'h00;
Memory[16022] = 8'h00;
Memory[16021] = 8'hCB;
Memory[16020] = 8'h20;
Memory[16027] = 8'h00;
Memory[16026] = 8'h00;
Memory[16025] = 8'hCC;
Memory[16024] = 8'h1A;
Memory[16031] = 8'h00;
Memory[16030] = 8'h00;
Memory[16029] = 8'hCE;
Memory[16028] = 8'h0E;
Memory[16035] = 8'h00;
Memory[16034] = 8'h00;
Memory[16033] = 8'hCF;
Memory[16032] = 8'h08;
Memory[16039] = 8'h00;
Memory[16038] = 8'h00;
Memory[16037] = 8'hD0;
Memory[16036] = 8'h02;
Memory[16043] = 8'h00;
Memory[16042] = 8'h00;
Memory[16041] = 8'hD0;
Memory[16040] = 8'hFC;
Memory[16047] = 8'h00;
Memory[16046] = 8'h00;
Memory[16045] = 8'hD1;
Memory[16044] = 8'hF6;
Memory[16051] = 8'h00;
Memory[16050] = 8'h00;
Memory[16049] = 8'hD2;
Memory[16048] = 8'hF0;
Memory[16055] = 8'h00;
Memory[16054] = 8'h00;
Memory[16053] = 8'hD3;
Memory[16052] = 8'hEA;
Memory[16059] = 8'h00;
Memory[16058] = 8'h00;
Memory[16057] = 8'hD4;
Memory[16056] = 8'hE4;
Memory[16063] = 8'h00;
Memory[16062] = 8'h00;
Memory[16061] = 8'hD5;
Memory[16060] = 8'hDE;
Memory[16067] = 8'h00;
Memory[16066] = 8'h00;
Memory[16065] = 8'hD6;
Memory[16064] = 8'hD8;
Memory[16071] = 8'h00;
Memory[16070] = 8'h00;
Memory[16069] = 8'hD7;
Memory[16068] = 8'hD2;
Memory[16075] = 8'h00;
Memory[16074] = 8'h00;
Memory[16073] = 8'hD8;
Memory[16072] = 8'hCC;
Memory[16079] = 8'h00;
Memory[16078] = 8'h00;
Memory[16077] = 8'hD9;
Memory[16076] = 8'hC6;
Memory[16083] = 8'h00;
Memory[16082] = 8'h00;
Memory[16081] = 8'hDA;
Memory[16080] = 8'hC0;
Memory[16087] = 8'h00;
Memory[16086] = 8'h00;
Memory[16085] = 8'hDC;
Memory[16084] = 8'hB4;
Memory[16091] = 8'h00;
Memory[16090] = 8'h00;
Memory[16089] = 8'hDE;
Memory[16088] = 8'hA8;
Memory[16095] = 8'h00;
Memory[16094] = 8'h00;
Memory[16093] = 8'hE2;
Memory[16092] = 8'h90;
Memory[16099] = 8'h00;
Memory[16098] = 8'h00;
Memory[16097] = 8'hE4;
Memory[16096] = 8'h84;
Memory[16103] = 8'h00;
Memory[16102] = 8'h00;
Memory[16101] = 8'hE6;
Memory[16100] = 8'h78;
Memory[16107] = 8'h00;
Memory[16106] = 8'h00;
Memory[16105] = 8'hEA;
Memory[16104] = 8'h60;
Memory[16111] = 8'h00;
Memory[16110] = 8'h00;
Memory[16109] = 8'hEE;
Memory[16108] = 8'h48;
Memory[16115] = 8'h00;
Memory[16114] = 8'h00;
Memory[16113] = 8'hF2;
Memory[16112] = 8'h30;
Memory[16119] = 8'h00;
Memory[16118] = 8'h00;
Memory[16117] = 8'hF6;
Memory[16116] = 8'h18;
Memory[16123] = 8'h00;
Memory[16122] = 8'h00;
Memory[16121] = 8'hFA;
Memory[16120] = 8'h00;
Memory[16127] = 8'h00;
Memory[16126] = 8'h00;
Memory[16125] = 8'hFB;
Memory[16124] = 8'hF4;
Memory[16131] = 8'h00;
Memory[16130] = 8'h00;
Memory[16129] = 8'hFD;
Memory[16128] = 8'hE8;
Memory[16135] = 8'h00;
Memory[16134] = 8'h01;
Memory[16133] = 8'h01;
Memory[16132] = 8'hD0;
Memory[16139] = 8'h00;
Memory[16138] = 8'h01;
Memory[16137] = 8'h03;
Memory[16136] = 8'hC4;
Memory[16143] = 8'h00;
Memory[16142] = 8'h01;
Memory[16141] = 8'h05;
Memory[16140] = 8'hB8;
Memory[16147] = 8'h00;
Memory[16146] = 8'h01;
Memory[16145] = 8'h13;
Memory[16144] = 8'h64;
Memory[16151] = 8'h00;
Memory[16150] = 8'h01;
Memory[16149] = 8'h15;
Memory[16148] = 8'h58;
Memory[16155] = 8'h00;
Memory[16154] = 8'h01;
Memory[16153] = 8'h17;
Memory[16152] = 8'h4C;
Memory[16159] = 8'h00;
Memory[16158] = 8'h01;
Memory[16157] = 8'h1A;
Memory[16156] = 8'h3A;
Memory[16163] = 8'h00;
Memory[16162] = 8'h01;
Memory[16161] = 8'h1A;
Memory[16160] = 8'hB7;
Memory[16167] = 8'h00;
Memory[16166] = 8'h01;
Memory[16165] = 8'h1B;
Memory[16164] = 8'h34;
Memory[16171] = 8'h00;
Memory[16170] = 8'h01;
Memory[16169] = 8'h1C;
Memory[16168] = 8'h2E;
Memory[16175] = 8'h00;
Memory[16174] = 8'h01;
Memory[16173] = 8'h1C;
Memory[16172] = 8'hAB;
Memory[16179] = 8'h00;
Memory[16178] = 8'h01;
Memory[16177] = 8'h1D;
Memory[16176] = 8'h28;
Memory[16183] = 8'h00;
Memory[16182] = 8'h01;
Memory[16181] = 8'h1D;
Memory[16180] = 8'hA5;
Memory[16187] = 8'h00;
Memory[16186] = 8'h01;
Memory[16185] = 8'h1E;
Memory[16184] = 8'h22;
Memory[16191] = 8'h00;
Memory[16190] = 8'h01;
Memory[16189] = 8'h1E;
Memory[16188] = 8'h9F;
Memory[16195] = 8'h00;
Memory[16194] = 8'h01;
Memory[16193] = 8'h1F;
Memory[16192] = 8'h1C;
Memory[16199] = 8'h00;
Memory[16198] = 8'h01;
Memory[16197] = 8'h1F;
Memory[16196] = 8'h99;
Memory[16203] = 8'h00;
Memory[16202] = 8'h01;
Memory[16201] = 8'h20;
Memory[16200] = 8'h16;
Memory[16207] = 8'h00;
Memory[16206] = 8'h01;
Memory[16205] = 8'h20;
Memory[16204] = 8'h93;
Memory[16211] = 8'h00;
Memory[16210] = 8'h01;
Memory[16209] = 8'h21;
Memory[16208] = 8'h10;
Memory[16215] = 8'h00;
Memory[16214] = 8'h01;
Memory[16213] = 8'h22;
Memory[16212] = 8'h0A;
Memory[16219] = 8'h00;
Memory[16218] = 8'h01;
Memory[16217] = 8'h22;
Memory[16216] = 8'h87;
Memory[16223] = 8'h00;
Memory[16222] = 8'h01;
Memory[16221] = 8'h23;
Memory[16220] = 8'h04;
Memory[16227] = 8'h00;
Memory[16226] = 8'h01;
Memory[16225] = 8'h23;
Memory[16224] = 8'hFE;
Memory[16231] = 8'h00;
Memory[16230] = 8'h01;
Memory[16229] = 8'h24;
Memory[16228] = 8'h7B;
Memory[16235] = 8'h00;
Memory[16234] = 8'h01;
Memory[16233] = 8'h24;
Memory[16232] = 8'hF8;
Memory[16239] = 8'h00;
Memory[16238] = 8'h01;
Memory[16237] = 8'h25;
Memory[16236] = 8'h75;
Memory[16243] = 8'h00;
Memory[16242] = 8'h01;
Memory[16241] = 8'h25;
Memory[16240] = 8'hF2;
Memory[16247] = 8'h00;
Memory[16246] = 8'h01;
Memory[16245] = 8'h26;
Memory[16244] = 8'h6F;
Memory[16251] = 8'h00;
Memory[16250] = 8'h01;
Memory[16249] = 8'h26;
Memory[16248] = 8'hEC;
Memory[16255] = 8'h00;
Memory[16254] = 8'h01;
Memory[16253] = 8'h27;
Memory[16252] = 8'h69;
Memory[16259] = 8'h00;
Memory[16258] = 8'h01;
Memory[16257] = 8'h27;
Memory[16256] = 8'hE6;
Memory[16263] = 8'h00;
Memory[16262] = 8'h01;
Memory[16261] = 8'h28;
Memory[16260] = 8'h63;
Memory[16267] = 8'h00;
Memory[16266] = 8'h01;
Memory[16265] = 8'h28;
Memory[16264] = 8'hE0;
Memory[16271] = 8'h00;
Memory[16270] = 8'h01;
Memory[16269] = 8'h29;
Memory[16268] = 8'hDA;
Memory[16275] = 8'h00;
Memory[16274] = 8'h01;
Memory[16273] = 8'h2A;
Memory[16272] = 8'h57;
Memory[16279] = 8'h00;
Memory[16278] = 8'h01;
Memory[16277] = 8'h2A;
Memory[16276] = 8'hD4;
Memory[16283] = 8'h00;
Memory[16282] = 8'h01;
Memory[16281] = 8'h2B;
Memory[16280] = 8'hCE;
Memory[16287] = 8'h00;
Memory[16286] = 8'h01;
Memory[16285] = 8'h2C;
Memory[16284] = 8'h4B;
Memory[16291] = 8'h00;
Memory[16290] = 8'h01;
Memory[16289] = 8'h2C;
Memory[16288] = 8'hC8;
Memory[16295] = 8'h00;
Memory[16294] = 8'h01;
Memory[16293] = 8'h2D;
Memory[16292] = 8'h45;
Memory[16299] = 8'h00;
Memory[16298] = 8'h01;
Memory[16297] = 8'h2D;
Memory[16296] = 8'hC2;
Memory[16303] = 8'h00;
Memory[16302] = 8'h01;
Memory[16301] = 8'h2E;
Memory[16300] = 8'h3F;
Memory[16307] = 8'h00;
Memory[16306] = 8'h01;
Memory[16305] = 8'h2E;
Memory[16304] = 8'hBC;
Memory[16311] = 8'h00;
Memory[16310] = 8'h01;
Memory[16309] = 8'h2F;
Memory[16308] = 8'h39;
Memory[16315] = 8'h00;
Memory[16314] = 8'h01;
Memory[16313] = 8'h2F;
Memory[16312] = 8'hB6;
Memory[16319] = 8'h00;
Memory[16318] = 8'h01;
Memory[16317] = 8'h30;
Memory[16316] = 8'h33;
Memory[16323] = 8'h00;
Memory[16322] = 8'h01;
Memory[16321] = 8'h30;
Memory[16320] = 8'hB0;
Memory[16327] = 8'h00;
Memory[16326] = 8'h01;
Memory[16325] = 8'h31;
Memory[16324] = 8'hAA;
Memory[16331] = 8'h00;
Memory[16330] = 8'h01;
Memory[16329] = 8'h32;
Memory[16328] = 8'h27;
Memory[16335] = 8'h00;
Memory[16334] = 8'h01;
Memory[16333] = 8'h32;
Memory[16332] = 8'hA4;
Memory[16339] = 8'h00;
Memory[16338] = 8'h01;
Memory[16337] = 8'h33;
Memory[16336] = 8'h9E;
Memory[16343] = 8'h00;
Memory[16342] = 8'h01;
Memory[16341] = 8'h34;
Memory[16340] = 8'h1B;
Memory[16347] = 8'h00;
Memory[16346] = 8'h01;
Memory[16345] = 8'h34;
Memory[16344] = 8'h98;
Memory[16351] = 8'h00;
Memory[16350] = 8'h01;
Memory[16349] = 8'h35;
Memory[16348] = 8'h15;
Memory[16355] = 8'h00;
Memory[16354] = 8'h01;
Memory[16353] = 8'h35;
Memory[16352] = 8'h92;
Memory[16359] = 8'h00;
Memory[16358] = 8'h01;
Memory[16357] = 8'h36;
Memory[16356] = 8'h0F;
Memory[16363] = 8'h00;
Memory[16362] = 8'h01;
Memory[16361] = 8'h36;
Memory[16360] = 8'h8C;
Memory[16367] = 8'h00;
Memory[16366] = 8'h01;
Memory[16365] = 8'h37;
Memory[16364] = 8'h09;
Memory[16371] = 8'h00;
Memory[16370] = 8'h01;
Memory[16369] = 8'h37;
Memory[16368] = 8'h86;
Memory[16375] = 8'h00;
Memory[16374] = 8'h01;
Memory[16373] = 8'h38;
Memory[16372] = 8'h03;
Memory[16379] = 8'h00;
Memory[16378] = 8'h01;
Memory[16377] = 8'h38;
Memory[16376] = 8'h80;
Memory[16383] = 8'h00;
Memory[16382] = 8'h01;
Memory[16381] = 8'h39;
Memory[16380] = 8'h7A;
Memory[16387] = 8'h00;
Memory[16386] = 8'h01;
Memory[16385] = 8'h39;
Memory[16384] = 8'hF7;
Memory[16391] = 8'h00;
Memory[16390] = 8'h01;
Memory[16389] = 8'h3A;
Memory[16388] = 8'h74;
Memory[16395] = 8'h00;
Memory[16394] = 8'h01;
Memory[16393] = 8'h3B;
Memory[16392] = 8'h6E;
Memory[16399] = 8'h00;
Memory[16398] = 8'h01;
Memory[16397] = 8'h3B;
Memory[16396] = 8'hEB;
Memory[16403] = 8'h00;
Memory[16402] = 8'h01;
Memory[16401] = 8'h3C;
Memory[16400] = 8'h68;
Memory[16407] = 8'h00;
Memory[16406] = 8'h01;
Memory[16405] = 8'h3C;
Memory[16404] = 8'hE5;
Memory[16411] = 8'h00;
Memory[16410] = 8'h01;
Memory[16409] = 8'h3D;
Memory[16408] = 8'h62;
Memory[16415] = 8'h00;
Memory[16414] = 8'h01;
Memory[16413] = 8'h3D;
Memory[16412] = 8'hDF;
Memory[16419] = 8'h00;
Memory[16418] = 8'h01;
Memory[16417] = 8'h3E;
Memory[16416] = 8'h5C;
Memory[16423] = 8'h00;
Memory[16422] = 8'h01;
Memory[16421] = 8'h3E;
Memory[16420] = 8'hD9;
Memory[16427] = 8'h00;
Memory[16426] = 8'h01;
Memory[16425] = 8'h3F;
Memory[16424] = 8'h56;
Memory[16431] = 8'h00;
Memory[16430] = 8'h01;
Memory[16429] = 8'h3F;
Memory[16428] = 8'hD3;
Memory[16435] = 8'h00;
Memory[16434] = 8'h01;
Memory[16433] = 8'h40;
Memory[16432] = 8'h50;
Memory[16439] = 8'h00;
Memory[16438] = 8'h01;
Memory[16437] = 8'h41;
Memory[16436] = 8'h4A;
Memory[16443] = 8'h00;
Memory[16442] = 8'h01;
Memory[16441] = 8'h41;
Memory[16440] = 8'hC7;
Memory[16447] = 8'h00;
Memory[16446] = 8'h01;
Memory[16445] = 8'h42;
Memory[16444] = 8'h44;
Memory[16451] = 8'h00;
Memory[16450] = 8'h01;
Memory[16449] = 8'h43;
Memory[16448] = 8'h3E;
Memory[16455] = 8'h00;
Memory[16454] = 8'h01;
Memory[16453] = 8'h43;
Memory[16452] = 8'hBB;
Memory[16459] = 8'h00;
Memory[16458] = 8'h01;
Memory[16457] = 8'h44;
Memory[16456] = 8'h38;
Memory[16463] = 8'h00;
Memory[16462] = 8'h01;
Memory[16461] = 8'h44;
Memory[16460] = 8'hB5;
Memory[16467] = 8'h00;
Memory[16466] = 8'h01;
Memory[16465] = 8'h45;
Memory[16464] = 8'h32;
Memory[16471] = 8'h00;
Memory[16470] = 8'h01;
Memory[16469] = 8'h45;
Memory[16468] = 8'hAF;
Memory[16475] = 8'h00;
Memory[16474] = 8'h01;
Memory[16473] = 8'h46;
Memory[16472] = 8'h2C;
Memory[16479] = 8'h00;
Memory[16478] = 8'h01;
Memory[16477] = 8'h46;
Memory[16476] = 8'hA9;
Memory[16483] = 8'h00;
Memory[16482] = 8'h01;
Memory[16481] = 8'h47;
Memory[16480] = 8'h26;
Memory[16487] = 8'h00;
Memory[16486] = 8'h01;
Memory[16485] = 8'h47;
Memory[16484] = 8'hA3;
Memory[16491] = 8'h00;
Memory[16490] = 8'h01;
Memory[16489] = 8'h48;
Memory[16488] = 8'h20;
Memory[16495] = 8'h00;
Memory[16494] = 8'h01;
Memory[16493] = 8'h49;
Memory[16492] = 8'h1A;
Memory[16499] = 8'h00;
Memory[16498] = 8'h01;
Memory[16497] = 8'h49;
Memory[16496] = 8'h97;
Memory[16503] = 8'h00;
Memory[16502] = 8'h01;
Memory[16501] = 8'h4A;
Memory[16500] = 8'h14;
Memory[16507] = 8'h00;
Memory[16506] = 8'h01;
Memory[16505] = 8'h4B;
Memory[16504] = 8'h0E;
Memory[16511] = 8'h00;
Memory[16510] = 8'h01;
Memory[16509] = 8'h4B;
Memory[16508] = 8'h8B;
Memory[16515] = 8'h00;
Memory[16514] = 8'h01;
Memory[16513] = 8'h4C;
Memory[16512] = 8'h08;
Memory[16519] = 8'h00;
Memory[16518] = 8'h01;
Memory[16517] = 8'h4C;
Memory[16516] = 8'h85;
Memory[16523] = 8'h00;
Memory[16522] = 8'h01;
Memory[16521] = 8'h4D;
Memory[16520] = 8'h02;
Memory[16527] = 8'h00;
Memory[16526] = 8'h01;
Memory[16525] = 8'h4D;
Memory[16524] = 8'h7F;
Memory[16531] = 8'h00;
Memory[16530] = 8'h01;
Memory[16529] = 8'h4D;
Memory[16528] = 8'hFC;
Memory[16535] = 8'h00;
Memory[16534] = 8'h01;
Memory[16533] = 8'h4E;
Memory[16532] = 8'h79;
Memory[16539] = 8'h00;
Memory[16538] = 8'h01;
Memory[16537] = 8'h4E;
Memory[16536] = 8'hF6;
Memory[16543] = 8'h00;
Memory[16542] = 8'h01;
Memory[16541] = 8'h4F;
Memory[16540] = 8'h73;
Memory[16547] = 8'h00;
Memory[16546] = 8'h01;
Memory[16545] = 8'h4F;
Memory[16544] = 8'hF0;
Memory[16551] = 8'h00;
Memory[16550] = 8'h01;
Memory[16549] = 8'h50;
Memory[16548] = 8'hEA;
Memory[16555] = 8'h00;
Memory[16554] = 8'h01;
Memory[16553] = 8'h51;
Memory[16552] = 8'h67;
Memory[16559] = 8'h00;
Memory[16558] = 8'h01;
Memory[16557] = 8'h51;
Memory[16556] = 8'hE4;
Memory[16563] = 8'h00;
Memory[16562] = 8'h01;
Memory[16561] = 8'h52;
Memory[16560] = 8'hDE;
Memory[16567] = 8'h00;
Memory[16566] = 8'h01;
Memory[16565] = 8'h53;
Memory[16564] = 8'h5B;
Memory[16571] = 8'h00;
Memory[16570] = 8'h01;
Memory[16569] = 8'h53;
Memory[16568] = 8'hD8;
Memory[16575] = 8'h00;
Memory[16574] = 8'h01;
Memory[16573] = 8'h54;
Memory[16572] = 8'h55;
Memory[16579] = 8'h00;
Memory[16578] = 8'h01;
Memory[16577] = 8'h54;
Memory[16576] = 8'hD2;
Memory[16583] = 8'h00;
Memory[16582] = 8'h01;
Memory[16581] = 8'h55;
Memory[16580] = 8'h4F;
Memory[16587] = 8'h00;
Memory[16586] = 8'h01;
Memory[16585] = 8'h55;
Memory[16584] = 8'hCC;
Memory[16591] = 8'h00;
Memory[16590] = 8'h01;
Memory[16589] = 8'h56;
Memory[16588] = 8'h49;
Memory[16595] = 8'h00;
Memory[16594] = 8'h01;
Memory[16593] = 8'h56;
Memory[16592] = 8'hC6;
Memory[16599] = 8'h00;
Memory[16598] = 8'h01;
Memory[16597] = 8'h57;
Memory[16596] = 8'h43;
Memory[16603] = 8'h00;
Memory[16602] = 8'h01;
Memory[16601] = 8'h57;
Memory[16600] = 8'hC0;
Memory[16607] = 8'h00;
Memory[16606] = 8'h01;
Memory[16605] = 8'h58;
Memory[16604] = 8'hBA;
Memory[16611] = 8'h00;
Memory[16610] = 8'h01;
Memory[16609] = 8'h59;
Memory[16608] = 8'h37;
Memory[16615] = 8'h00;
Memory[16614] = 8'h01;
Memory[16613] = 8'h59;
Memory[16612] = 8'hB4;
Memory[16619] = 8'h00;
Memory[16618] = 8'h01;
Memory[16617] = 8'h5A;
Memory[16616] = 8'hAE;
Memory[16623] = 8'h00;
Memory[16622] = 8'h01;
Memory[16621] = 8'h5B;
Memory[16620] = 8'h2B;
Memory[16627] = 8'h00;
Memory[16626] = 8'h01;
Memory[16625] = 8'h5B;
Memory[16624] = 8'hA8;
Memory[16631] = 8'h00;
Memory[16630] = 8'h01;
Memory[16629] = 8'h5C;
Memory[16628] = 8'h25;
Memory[16635] = 8'h00;
Memory[16634] = 8'h01;
Memory[16633] = 8'h5C;
Memory[16632] = 8'hA2;
Memory[16639] = 8'h00;
Memory[16638] = 8'h01;
Memory[16637] = 8'h5D;
Memory[16636] = 8'h1F;
Memory[16643] = 8'h00;
Memory[16642] = 8'h01;
Memory[16641] = 8'h5D;
Memory[16640] = 8'h9C;
Memory[16647] = 8'h00;
Memory[16646] = 8'h01;
Memory[16645] = 8'h5E;
Memory[16644] = 8'h19;
Memory[16651] = 8'h00;
Memory[16650] = 8'h01;
Memory[16649] = 8'h5E;
Memory[16648] = 8'h96;
Memory[16655] = 8'h00;
Memory[16654] = 8'h01;
Memory[16653] = 8'h5F;
Memory[16652] = 8'h13;
Memory[16659] = 8'h00;
Memory[16658] = 8'h01;
Memory[16657] = 8'h5F;
Memory[16656] = 8'h90;
Memory[16663] = 8'h00;
Memory[16662] = 8'h01;
Memory[16661] = 8'h60;
Memory[16660] = 8'h8A;
Memory[16667] = 8'h00;
Memory[16666] = 8'h01;
Memory[16665] = 8'h61;
Memory[16664] = 8'h07;
Memory[16671] = 8'h00;
Memory[16670] = 8'h01;
Memory[16669] = 8'h61;
Memory[16668] = 8'h84;
Memory[16675] = 8'h00;
Memory[16674] = 8'h01;
Memory[16673] = 8'h62;
Memory[16672] = 8'h7E;
Memory[16679] = 8'h00;
Memory[16678] = 8'h01;
Memory[16677] = 8'h62;
Memory[16676] = 8'hFB;
Memory[16683] = 8'h00;
Memory[16682] = 8'h01;
Memory[16681] = 8'h63;
Memory[16680] = 8'h78;
Memory[16687] = 8'h00;
Memory[16686] = 8'h01;
Memory[16685] = 8'h63;
Memory[16684] = 8'hF5;
Memory[16691] = 8'h00;
Memory[16690] = 8'h01;
Memory[16689] = 8'h64;
Memory[16688] = 8'h72;
Memory[16695] = 8'h00;
Memory[16694] = 8'h01;
Memory[16693] = 8'h64;
Memory[16692] = 8'hEF;
Memory[16699] = 8'h00;
Memory[16698] = 8'h01;
Memory[16697] = 8'h65;
Memory[16696] = 8'h6C;
Memory[16703] = 8'h00;
Memory[16702] = 8'h01;
Memory[16701] = 8'h65;
Memory[16700] = 8'hE9;
Memory[16707] = 8'h00;
Memory[16706] = 8'h01;
Memory[16705] = 8'h66;
Memory[16704] = 8'h66;
Memory[16711] = 8'h00;
Memory[16710] = 8'h01;
Memory[16709] = 8'h66;
Memory[16708] = 8'hE3;
Memory[16715] = 8'h00;
Memory[16714] = 8'h01;
Memory[16713] = 8'h67;
Memory[16712] = 8'h60;
Memory[16719] = 8'h00;
Memory[16718] = 8'h01;
Memory[16717] = 8'h68;
Memory[16716] = 8'h5A;
Memory[16723] = 8'h00;
Memory[16722] = 8'h01;
Memory[16721] = 8'h68;
Memory[16720] = 8'hD7;
Memory[16727] = 8'h00;
Memory[16726] = 8'h01;
Memory[16725] = 8'h69;
Memory[16724] = 8'h54;
Memory[16731] = 8'h00;
Memory[16730] = 8'h01;
Memory[16729] = 8'h6A;
Memory[16728] = 8'h4E;
Memory[16735] = 8'h00;
Memory[16734] = 8'h01;
Memory[16733] = 8'h6A;
Memory[16732] = 8'hCB;
Memory[16739] = 8'h00;
Memory[16738] = 8'h01;
Memory[16737] = 8'h6B;
Memory[16736] = 8'h48;
Memory[16743] = 8'h00;
Memory[16742] = 8'h01;
Memory[16741] = 8'h6B;
Memory[16740] = 8'hC5;
Memory[16747] = 8'h00;
Memory[16746] = 8'h01;
Memory[16745] = 8'h6C;
Memory[16744] = 8'h42;
Memory[16751] = 8'h00;
Memory[16750] = 8'h01;
Memory[16749] = 8'h6C;
Memory[16748] = 8'hBF;
Memory[16755] = 8'h00;
Memory[16754] = 8'h01;
Memory[16753] = 8'h6D;
Memory[16752] = 8'h3C;
Memory[16759] = 8'h00;
Memory[16758] = 8'h01;
Memory[16757] = 8'h6D;
Memory[16756] = 8'hB9;
Memory[16763] = 8'h00;
Memory[16762] = 8'h01;
Memory[16761] = 8'h6E;
Memory[16760] = 8'h36;
Memory[16767] = 8'h00;
Memory[16766] = 8'h01;
Memory[16765] = 8'h6E;
Memory[16764] = 8'hB3;
Memory[16771] = 8'h00;
Memory[16770] = 8'h01;
Memory[16769] = 8'h6F;
Memory[16768] = 8'h30;
Memory[16775] = 8'h00;
Memory[16774] = 8'h01;
Memory[16773] = 8'h70;
Memory[16772] = 8'h2A;
Memory[16779] = 8'h00;
Memory[16778] = 8'h01;
Memory[16777] = 8'h70;
Memory[16776] = 8'hA7;
Memory[16783] = 8'h00;
Memory[16782] = 8'h01;
Memory[16781] = 8'h71;
Memory[16780] = 8'h24;
Memory[16787] = 8'h00;
Memory[16786] = 8'h01;
Memory[16785] = 8'h72;
Memory[16784] = 8'h1E;
Memory[16791] = 8'h00;
Memory[16790] = 8'h01;
Memory[16789] = 8'h72;
Memory[16788] = 8'h9B;
Memory[16795] = 8'h00;
Memory[16794] = 8'h01;
Memory[16793] = 8'h73;
Memory[16792] = 8'h18;
Memory[16799] = 8'h00;
Memory[16798] = 8'h01;
Memory[16797] = 8'h73;
Memory[16796] = 8'h95;
Memory[16803] = 8'h00;
Memory[16802] = 8'h01;
Memory[16801] = 8'h74;
Memory[16800] = 8'h12;
Memory[16807] = 8'h00;
Memory[16806] = 8'h01;
Memory[16805] = 8'h74;
Memory[16804] = 8'h8F;
Memory[16811] = 8'h00;
Memory[16810] = 8'h01;
Memory[16809] = 8'h75;
Memory[16808] = 8'h0C;
Memory[16815] = 8'h00;
Memory[16814] = 8'h01;
Memory[16813] = 8'h75;
Memory[16812] = 8'h89;
Memory[16819] = 8'h00;
Memory[16818] = 8'h01;
Memory[16817] = 8'h76;
Memory[16816] = 8'h06;
Memory[16823] = 8'h00;
Memory[16822] = 8'h01;
Memory[16821] = 8'h76;
Memory[16820] = 8'h83;
Memory[16827] = 8'h00;
Memory[16826] = 8'h01;
Memory[16825] = 8'h77;
Memory[16824] = 8'h00;
Memory[16831] = 8'h00;
Memory[16830] = 8'h01;
Memory[16829] = 8'h77;
Memory[16828] = 8'hFA;
Memory[16835] = 8'h00;
Memory[16834] = 8'h01;
Memory[16833] = 8'h78;
Memory[16832] = 8'h77;
Memory[16839] = 8'h00;
Memory[16838] = 8'h01;
Memory[16837] = 8'h78;
Memory[16836] = 8'hF4;
Memory[16843] = 8'h00;
Memory[16842] = 8'h01;
Memory[16841] = 8'h79;
Memory[16840] = 8'hEE;
Memory[16847] = 8'h00;
Memory[16846] = 8'h01;
Memory[16845] = 8'h7A;
Memory[16844] = 8'h6B;
Memory[16851] = 8'h00;
Memory[16850] = 8'h01;
Memory[16849] = 8'h7A;
Memory[16848] = 8'hE8;
Memory[16855] = 8'h00;
Memory[16854] = 8'h01;
Memory[16853] = 8'h7B;
Memory[16852] = 8'h65;
Memory[16859] = 8'h00;
Memory[16858] = 8'h01;
Memory[16857] = 8'h7B;
Memory[16856] = 8'hE2;
Memory[16863] = 8'h00;
Memory[16862] = 8'h01;
Memory[16861] = 8'h7C;
Memory[16860] = 8'h5F;
Memory[16867] = 8'h00;
Memory[16866] = 8'h01;
Memory[16865] = 8'h7C;
Memory[16864] = 8'hDC;
Memory[16871] = 8'h00;
Memory[16870] = 8'h01;
Memory[16869] = 8'h7D;
Memory[16868] = 8'h59;
Memory[16875] = 8'h00;
Memory[16874] = 8'h01;
Memory[16873] = 8'h7D;
Memory[16872] = 8'hD6;
Memory[16879] = 8'h00;
Memory[16878] = 8'h01;
Memory[16877] = 8'h7E;
Memory[16876] = 8'h53;
Memory[16883] = 8'h00;
Memory[16882] = 8'h01;
Memory[16881] = 8'h7E;
Memory[16880] = 8'hD0;
Memory[16887] = 8'h00;
Memory[16886] = 8'h01;
Memory[16885] = 8'h7F;
Memory[16884] = 8'hCA;
Memory[16891] = 8'h00;
Memory[16890] = 8'h01;
Memory[16889] = 8'h80;
Memory[16888] = 8'h47;
Memory[16895] = 8'h00;
Memory[16894] = 8'h01;
Memory[16893] = 8'h80;
Memory[16892] = 8'hC4;
Memory[16899] = 8'h00;
Memory[16898] = 8'h01;
Memory[16897] = 8'h81;
Memory[16896] = 8'hBE;
Memory[16903] = 8'h00;
Memory[16902] = 8'h01;
Memory[16901] = 8'h82;
Memory[16900] = 8'h3B;
Memory[16907] = 8'h00;
Memory[16906] = 8'h01;
Memory[16905] = 8'h82;
Memory[16904] = 8'hB8;
Memory[16911] = 8'h00;
Memory[16910] = 8'h01;
Memory[16909] = 8'h83;
Memory[16908] = 8'h35;
Memory[16915] = 8'h00;
Memory[16914] = 8'h01;
Memory[16913] = 8'h83;
Memory[16912] = 8'hB2;
Memory[16919] = 8'h00;
Memory[16918] = 8'h01;
Memory[16917] = 8'h84;
Memory[16916] = 8'h2F;
Memory[16923] = 8'h00;
Memory[16922] = 8'h01;
Memory[16921] = 8'h84;
Memory[16920] = 8'hAC;
Memory[16927] = 8'h00;
Memory[16926] = 8'h01;
Memory[16925] = 8'h85;
Memory[16924] = 8'h29;
Memory[16931] = 8'h00;
Memory[16930] = 8'h01;
Memory[16929] = 8'h85;
Memory[16928] = 8'hA6;
Memory[16935] = 8'h00;
Memory[16934] = 8'h01;
Memory[16933] = 8'h86;
Memory[16932] = 8'h23;
Memory[16939] = 8'h00;
Memory[16938] = 8'h01;
Memory[16937] = 8'h86;
Memory[16936] = 8'hA0;
Memory[16943] = 8'h00;
Memory[16942] = 8'h01;
Memory[16941] = 8'h87;
Memory[16940] = 8'h9A;
Memory[16947] = 8'h00;
Memory[16946] = 8'h01;
Memory[16945] = 8'h88;
Memory[16944] = 8'h17;
Memory[16951] = 8'h00;
Memory[16950] = 8'h01;
Memory[16949] = 8'h88;
Memory[16948] = 8'h94;
Memory[16955] = 8'h00;
Memory[16954] = 8'h01;
Memory[16953] = 8'h89;
Memory[16952] = 8'h8E;
Memory[16959] = 8'h00;
Memory[16958] = 8'h01;
Memory[16957] = 8'h8A;
Memory[16956] = 8'h0B;
Memory[16963] = 8'h00;
Memory[16962] = 8'h01;
Memory[16961] = 8'h8A;
Memory[16960] = 8'h88;
Memory[16967] = 8'h00;
Memory[16966] = 8'h01;
Memory[16965] = 8'h8B;
Memory[16964] = 8'h05;
Memory[16971] = 8'h00;
Memory[16970] = 8'h01;
Memory[16969] = 8'h8B;
Memory[16968] = 8'h82;
Memory[16975] = 8'h00;
Memory[16974] = 8'h01;
Memory[16973] = 8'h8B;
Memory[16972] = 8'hFF;
Memory[16979] = 8'h00;
Memory[16978] = 8'h01;
Memory[16977] = 8'h8C;
Memory[16976] = 8'h7C;
Memory[16983] = 8'h00;
Memory[16982] = 8'h01;
Memory[16981] = 8'h8C;
Memory[16980] = 8'hF9;
Memory[16987] = 8'h00;
Memory[16986] = 8'h01;
Memory[16985] = 8'h8D;
Memory[16984] = 8'h76;
Memory[16991] = 8'h00;
Memory[16990] = 8'h01;
Memory[16989] = 8'h8D;
Memory[16988] = 8'hF3;
Memory[16995] = 8'h00;
Memory[16994] = 8'h01;
Memory[16993] = 8'h8E;
Memory[16992] = 8'h70;
Memory[16999] = 8'h00;
Memory[16998] = 8'h01;
Memory[16997] = 8'h8F;
Memory[16996] = 8'h6A;
Memory[17003] = 8'h00;
Memory[17002] = 8'h01;
Memory[17001] = 8'h8F;
Memory[17000] = 8'hE7;
Memory[17007] = 8'h00;
Memory[17006] = 8'h01;
Memory[17005] = 8'h90;
Memory[17004] = 8'h64;
Memory[17011] = 8'h00;
Memory[17010] = 8'h01;
Memory[17009] = 8'h91;
Memory[17008] = 8'h5E;
Memory[17015] = 8'h00;
Memory[17014] = 8'h01;
Memory[17013] = 8'h91;
Memory[17012] = 8'hDB;
Memory[17019] = 8'h00;
Memory[17018] = 8'h01;
Memory[17017] = 8'h92;
Memory[17016] = 8'h58;
Memory[17023] = 8'h00;
Memory[17022] = 8'h01;
Memory[17021] = 8'h92;
Memory[17020] = 8'hD5;
Memory[17027] = 8'h00;
Memory[17026] = 8'h01;
Memory[17025] = 8'h93;
Memory[17024] = 8'h52;
Memory[17031] = 8'h00;
Memory[17030] = 8'h01;
Memory[17029] = 8'h93;
Memory[17028] = 8'hCF;
Memory[17035] = 8'h00;
Memory[17034] = 8'h01;
Memory[17033] = 8'h94;
Memory[17032] = 8'h4C;
Memory[17039] = 8'h00;
Memory[17038] = 8'h01;
Memory[17037] = 8'h94;
Memory[17036] = 8'hC9;
Memory[17043] = 8'h00;
Memory[17042] = 8'h01;
Memory[17041] = 8'h95;
Memory[17040] = 8'h46;
Memory[17047] = 8'h00;
Memory[17046] = 8'h01;
Memory[17045] = 8'h95;
Memory[17044] = 8'hC3;
Memory[17051] = 8'h00;
Memory[17050] = 8'h01;
Memory[17049] = 8'h96;
Memory[17048] = 8'h40;
Memory[17055] = 8'h00;
Memory[17054] = 8'h01;
Memory[17053] = 8'h99;
Memory[17052] = 8'h2E;
Memory[17059] = 8'h00;
Memory[17058] = 8'h01;
Memory[17057] = 8'h9B;
Memory[17056] = 8'h22;
Memory[17063] = 8'h00;
Memory[17062] = 8'h01;
Memory[17061] = 8'h9C;
Memory[17060] = 8'h1C;
Memory[17067] = 8'h00;
Memory[17066] = 8'h01;
Memory[17065] = 8'h9D;
Memory[17064] = 8'h16;
Memory[17071] = 8'h00;
Memory[17070] = 8'h01;
Memory[17069] = 8'h9E;
Memory[17068] = 8'h10;
Memory[17075] = 8'h00;
Memory[17074] = 8'h01;
Memory[17073] = 8'hA2;
Memory[17072] = 8'hF2;
Memory[17079] = 8'h00;
Memory[17078] = 8'h01;
Memory[17077] = 8'hA3;
Memory[17076] = 8'hEC;
Memory[17083] = 8'h00;
Memory[17082] = 8'h01;
Memory[17081] = 8'hA4;
Memory[17080] = 8'hE6;
Memory[17087] = 8'h00;
Memory[17086] = 8'h01;
Memory[17085] = 8'hA5;
Memory[17084] = 8'hE0;
Memory[17091] = 8'h00;
Memory[17090] = 8'h01;
Memory[17089] = 8'hA9;
Memory[17088] = 8'hC8;
Memory[17095] = 8'h00;
Memory[17094] = 8'h01;
Memory[17093] = 8'hAE;
Memory[17092] = 8'hAA;
Memory[17099] = 8'h00;
Memory[17098] = 8'h01;
Memory[17097] = 8'hAF;
Memory[17096] = 8'hA4;
Memory[17103] = 8'h00;
Memory[17102] = 8'h01;
Memory[17101] = 8'hB0;
Memory[17100] = 8'h9E;
Memory[17107] = 8'h00;
Memory[17106] = 8'h01;
Memory[17105] = 8'hB1;
Memory[17104] = 8'h98;
Memory[17111] = 8'h00;
Memory[17110] = 8'h01;
Memory[17109] = 8'hB8;
Memory[17108] = 8'h6E;
Memory[17115] = 8'h00;
Memory[17114] = 8'h01;
Memory[17113] = 8'hBA;
Memory[17112] = 8'h62;
Memory[17119] = 8'h00;
Memory[17118] = 8'h01;
Memory[17117] = 8'hBB;
Memory[17116] = 8'h5C;
Memory[17123] = 8'h00;
Memory[17122] = 8'h01;
Memory[17121] = 8'hBC;
Memory[17120] = 8'h56;
Memory[17127] = 8'h00;
Memory[17126] = 8'h01;
Memory[17125] = 8'hBD;
Memory[17124] = 8'h50;
Memory[17131] = 8'h00;
Memory[17130] = 8'h01;
Memory[17129] = 8'hC2;
Memory[17128] = 8'h32;
Memory[17135] = 8'h00;
Memory[17134] = 8'h01;
Memory[17133] = 8'hC3;
Memory[17132] = 8'h2C;
Memory[17139] = 8'h00;
Memory[17138] = 8'h01;
Memory[17137] = 8'hC4;
Memory[17136] = 8'h26;
Memory[17143] = 8'h00;
Memory[17142] = 8'h01;
Memory[17141] = 8'hC5;
Memory[17140] = 8'h20;
Memory[17147] = 8'h00;
Memory[17146] = 8'h01;
Memory[17145] = 8'hC6;
Memory[17144] = 8'h1A;
Memory[17151] = 8'h00;
Memory[17150] = 8'h01;
Memory[17149] = 8'hC7;
Memory[17148] = 8'h14;
Memory[17155] = 8'h00;
Memory[17154] = 8'h01;
Memory[17153] = 8'hC8;
Memory[17152] = 8'h0E;
Memory[17159] = 8'h00;
Memory[17158] = 8'h01;
Memory[17157] = 8'hC9;
Memory[17156] = 8'h08;
Memory[17163] = 8'h00;
Memory[17162] = 8'h01;
Memory[17161] = 8'hCC;
Memory[17160] = 8'hF0;
Memory[17167] = 8'h00;
Memory[17166] = 8'h01;
Memory[17165] = 8'hCE;
Memory[17164] = 8'hE4;
Memory[17171] = 8'h00;
Memory[17170] = 8'h01;
Memory[17169] = 8'hD0;
Memory[17168] = 8'hD8;
Memory[17175] = 8'h00;
Memory[17174] = 8'h01;
Memory[17173] = 8'hD4;
Memory[17172] = 8'hC0;
Memory[17179] = 8'h00;
Memory[17178] = 8'h01;
Memory[17177] = 8'hD7;
Memory[17176] = 8'hAE;
Memory[17183] = 8'h00;
Memory[17182] = 8'h01;
Memory[17181] = 8'hD9;
Memory[17180] = 8'hA2;
Memory[17187] = 8'h00;
Memory[17186] = 8'h01;
Memory[17185] = 8'hDA;
Memory[17184] = 8'h9C;
Memory[17191] = 8'h00;
Memory[17190] = 8'h01;
Memory[17189] = 8'hDB;
Memory[17188] = 8'h96;
Memory[17195] = 8'h00;
Memory[17194] = 8'h01;
Memory[17193] = 8'hDC;
Memory[17192] = 8'h90;
Memory[17199] = 8'h00;
Memory[17198] = 8'h01;
Memory[17197] = 8'hE1;
Memory[17196] = 8'h72;
Memory[17203] = 8'h00;
Memory[17202] = 8'h01;
Memory[17201] = 8'hE2;
Memory[17200] = 8'h6C;
Memory[17207] = 8'h00;
Memory[17206] = 8'h01;
Memory[17205] = 8'hE3;
Memory[17204] = 8'h66;
Memory[17211] = 8'h00;
Memory[17210] = 8'h01;
Memory[17209] = 8'hE4;
Memory[17208] = 8'h60;
Memory[17215] = 8'h00;
Memory[17214] = 8'h01;
Memory[17213] = 8'hE8;
Memory[17212] = 8'h48;
Memory[17219] = 8'h00;
Memory[17218] = 8'h01;
Memory[17217] = 8'hED;
Memory[17216] = 8'h2A;
Memory[17223] = 8'h00;
Memory[17222] = 8'h01;
Memory[17221] = 8'hEE;
Memory[17220] = 8'h24;
Memory[17227] = 8'h00;
Memory[17226] = 8'h01;
Memory[17225] = 8'hEF;
Memory[17224] = 8'h1E;
Memory[17231] = 8'h00;
Memory[17230] = 8'h01;
Memory[17229] = 8'hF0;
Memory[17228] = 8'h18;
Memory[17235] = 8'h00;
Memory[17234] = 8'h01;
Memory[17233] = 8'hF6;
Memory[17232] = 8'hEE;
Memory[17239] = 8'h00;
Memory[17238] = 8'h01;
Memory[17237] = 8'hF8;
Memory[17236] = 8'hE2;
Memory[17243] = 8'h00;
Memory[17242] = 8'h01;
Memory[17241] = 8'hF9;
Memory[17240] = 8'hDC;
Memory[17247] = 8'h00;
Memory[17246] = 8'h01;
Memory[17245] = 8'hFA;
Memory[17244] = 8'hD6;
Memory[17251] = 8'h00;
Memory[17250] = 8'h01;
Memory[17249] = 8'hFB;
Memory[17248] = 8'hD0;
Memory[17255] = 8'h00;
Memory[17254] = 8'h02;
Memory[17253] = 8'h00;
Memory[17252] = 8'hB2;
Memory[17259] = 8'h00;
Memory[17258] = 8'h02;
Memory[17257] = 8'h01;
Memory[17256] = 8'hAC;
Memory[17263] = 8'h00;
Memory[17262] = 8'h02;
Memory[17261] = 8'h02;
Memory[17260] = 8'hA6;
Memory[17267] = 8'h00;
Memory[17266] = 8'h02;
Memory[17265] = 8'h03;
Memory[17264] = 8'hA0;
Memory[17271] = 8'h00;
Memory[17270] = 8'h02;
Memory[17269] = 8'h04;
Memory[17268] = 8'h9A;
Memory[17275] = 8'h00;
Memory[17274] = 8'h02;
Memory[17273] = 8'h05;
Memory[17272] = 8'h94;
Memory[17279] = 8'h00;
Memory[17278] = 8'h02;
Memory[17277] = 8'h06;
Memory[17276] = 8'h8E;
Memory[17283] = 8'h00;
Memory[17282] = 8'h02;
Memory[17281] = 8'h07;
Memory[17280] = 8'h88;
Memory[17287] = 8'h00;
Memory[17286] = 8'h02;
Memory[17285] = 8'h0B;
Memory[17284] = 8'h70;
Memory[17291] = 8'h00;
Memory[17290] = 8'h02;
Memory[17289] = 8'h0D;
Memory[17288] = 8'h64;
Memory[17295] = 8'h00;
Memory[17294] = 8'h02;
Memory[17293] = 8'h0F;
Memory[17292] = 8'h58;
Memory[17299] = 8'h00;
Memory[17298] = 8'h02;
Memory[17297] = 8'h13;
Memory[17296] = 8'h40;
Memory[17303] = 8'h00;
Memory[17302] = 8'h02;
Memory[17301] = 8'h17;
Memory[17300] = 8'h28;
Memory[17307] = 8'h00;
Memory[17306] = 8'h02;
Memory[17305] = 8'h1B;
Memory[17304] = 8'h10;
Memory[17311] = 8'h00;
Memory[17310] = 8'h02;
Memory[17309] = 8'h1E;
Memory[17308] = 8'hF8;
Memory[17315] = 8'h00;
Memory[17314] = 8'h02;
Memory[17313] = 8'h22;
Memory[17312] = 8'hE0;
Memory[17319] = 8'h00;
Memory[17318] = 8'h02;
Memory[17317] = 8'h26;
Memory[17316] = 8'hC8;
Memory[17323] = 8'h00;
Memory[17322] = 8'h02;
Memory[17321] = 8'h2A;
Memory[17320] = 8'hB0;
Memory[17327] = 8'h00;
Memory[17326] = 8'h02;
Memory[17325] = 8'h2E;
Memory[17324] = 8'h98;
Memory[17331] = 8'h00;
Memory[17330] = 8'h02;
Memory[17329] = 8'h32;
Memory[17328] = 8'h80;
Memory[17335] = 8'h00;
Memory[17334] = 8'h02;
Memory[17333] = 8'h36;
Memory[17332] = 8'h68;
Memory[17339] = 8'h00;
Memory[17338] = 8'h02;
Memory[17337] = 8'h3A;
Memory[17336] = 8'h50;
Memory[17343] = 8'h00;
Memory[17342] = 8'h02;
Memory[17341] = 8'h3E;
Memory[17340] = 8'h38;
Memory[17347] = 8'h00;
Memory[17346] = 8'h02;
Memory[17345] = 8'h42;
Memory[17344] = 8'h20;
Memory[17351] = 8'h00;
Memory[17350] = 8'h02;
Memory[17349] = 8'h44;
Memory[17348] = 8'h14;
Memory[17355] = 8'h00;
Memory[17354] = 8'h02;
Memory[17353] = 8'h46;
Memory[17352] = 8'h08;
Memory[17359] = 8'h00;
Memory[17358] = 8'h02;
Memory[17357] = 8'h47;
Memory[17356] = 8'hFC;
Memory[17363] = 8'h00;
Memory[17362] = 8'h02;
Memory[17361] = 8'h49;
Memory[17360] = 8'hF0;
Memory[17367] = 8'h00;
Memory[17366] = 8'h02;
Memory[17365] = 8'h4D;
Memory[17364] = 8'hD8;
Memory[17371] = 8'h00;
Memory[17370] = 8'h02;
Memory[17369] = 8'h51;
Memory[17368] = 8'hC0;
Memory[17375] = 8'h00;
Memory[17374] = 8'h02;
Memory[17373] = 8'h59;
Memory[17372] = 8'h90;
Memory[17379] = 8'h00;
Memory[17378] = 8'h00;
Memory[17377] = 8'h01;
Memory[17376] = 8'h25;
Memory[17383] = 8'h00;
Memory[17382] = 8'h00;
Memory[17381] = 8'h00;
Memory[17380] = 8'hDC;
Memory[17387] = 8'h00;
Memory[17386] = 8'h00;
Memory[17385] = 8'h00;
Memory[17384] = 8'hF6;
Memory[17391] = 8'h00;
Memory[17390] = 8'h00;
Memory[17389] = 8'h00;
Memory[17388] = 8'hB8;
Memory[17395] = 8'h00;
Memory[17394] = 8'h00;
Memory[17393] = 8'h00;
Memory[17392] = 8'hC3;
Memory[17399] = 8'h00;
Memory[17398] = 8'h00;
Memory[17397] = 8'h00;
Memory[17396] = 8'h92;
Memory[17403] = 8'h00;
Memory[17402] = 8'h00;
Memory[17401] = 8'h00;
Memory[17400] = 8'hC3;
Memory[17407] = 8'h00;
Memory[17406] = 8'h00;
Memory[17405] = 8'h00;
Memory[17404] = 8'hDC;
Memory[17411] = 8'h00;
Memory[17410] = 8'h00;
Memory[17409] = 8'h01;
Memory[17408] = 8'h71;
Memory[17415] = 8'h00;
Memory[17414] = 8'h00;
Memory[17413] = 8'h01;
Memory[17412] = 8'h49;
Memory[17419] = 8'h00;
Memory[17418] = 8'h00;
Memory[17417] = 8'h01;
Memory[17416] = 8'h25;
Memory[17423] = 8'h00;
Memory[17422] = 8'h00;
Memory[17421] = 8'h01;
Memory[17420] = 8'h15;
Memory[17427] = 8'h00;
Memory[17426] = 8'h00;
Memory[17425] = 8'h00;
Memory[17424] = 8'hF6;
Memory[17431] = 8'h00;
Memory[17430] = 8'h00;
Memory[17429] = 8'h00;
Memory[17428] = 8'hDC;
Memory[17435] = 8'h00;
Memory[17434] = 8'h00;
Memory[17433] = 8'h00;
Memory[17432] = 8'hF6;
Memory[17439] = 8'h00;
Memory[17438] = 8'h00;
Memory[17437] = 8'h01;
Memory[17436] = 8'h15;
Memory[17443] = 8'h00;
Memory[17442] = 8'h00;
Memory[17441] = 8'h01;
Memory[17440] = 8'h25;
Memory[17447] = 8'h00;
Memory[17446] = 8'h00;
Memory[17445] = 8'h01;
Memory[17444] = 8'h15;
Memory[17451] = 8'h00;
Memory[17450] = 8'h00;
Memory[17449] = 8'h00;
Memory[17448] = 8'hF6;
Memory[17455] = 8'h00;
Memory[17454] = 8'h00;
Memory[17453] = 8'h00;
Memory[17452] = 8'hDC;
Memory[17459] = 8'h00;
Memory[17458] = 8'h00;
Memory[17457] = 8'h00;
Memory[17456] = 8'hC3;
Memory[17463] = 8'h00;
Memory[17462] = 8'h00;
Memory[17461] = 8'h00;
Memory[17460] = 8'hB8;
Memory[17467] = 8'h00;
Memory[17466] = 8'h00;
Memory[17465] = 8'h00;
Memory[17464] = 8'hC3;
Memory[17471] = 8'h00;
Memory[17470] = 8'h00;
Memory[17469] = 8'h00;
Memory[17468] = 8'hA4;
Memory[17475] = 8'h00;
Memory[17474] = 8'h00;
Memory[17473] = 8'h00;
Memory[17472] = 8'h92;
Memory[17479] = 8'h00;
Memory[17478] = 8'h00;
Memory[17477] = 8'h00;
Memory[17476] = 8'hB8;
Memory[17483] = 8'h00;
Memory[17482] = 8'h00;
Memory[17481] = 8'h00;
Memory[17480] = 8'hDC;
Memory[17487] = 8'h00;
Memory[17486] = 8'h00;
Memory[17485] = 8'h00;
Memory[17484] = 8'hC3;
Memory[17491] = 8'h00;
Memory[17490] = 8'h00;
Memory[17489] = 8'h00;
Memory[17488] = 8'hB8;
Memory[17495] = 8'h00;
Memory[17494] = 8'h00;
Memory[17493] = 8'h00;
Memory[17492] = 8'h92;
Memory[17499] = 8'h00;
Memory[17498] = 8'h00;
Memory[17497] = 8'h00;
Memory[17496] = 8'hB8;
Memory[17503] = 8'h00;
Memory[17502] = 8'h00;
Memory[17501] = 8'h00;
Memory[17500] = 8'hA4;
Memory[17507] = 8'h00;
Memory[17506] = 8'h00;
Memory[17505] = 8'h00;
Memory[17504] = 8'h92;
Memory[17511] = 8'h00;
Memory[17510] = 8'h00;
Memory[17509] = 8'h00;
Memory[17508] = 8'hF6;
Memory[17515] = 8'h00;
Memory[17514] = 8'h00;
Memory[17513] = 8'h00;
Memory[17512] = 8'h92;
Memory[17519] = 8'h00;
Memory[17518] = 8'h00;
Memory[17517] = 8'h00;
Memory[17516] = 8'hDC;
Memory[17523] = 8'h00;
Memory[17522] = 8'h00;
Memory[17521] = 8'h00;
Memory[17520] = 8'hC3;
Memory[17527] = 8'h00;
Memory[17526] = 8'h00;
Memory[17525] = 8'h00;
Memory[17524] = 8'hF6;
Memory[17531] = 8'h00;
Memory[17530] = 8'h00;
Memory[17529] = 8'h00;
Memory[17528] = 8'hDC;
Memory[17535] = 8'h00;
Memory[17534] = 8'h00;
Memory[17533] = 8'h00;
Memory[17532] = 8'hC3;
Memory[17539] = 8'h00;
Memory[17538] = 8'h00;
Memory[17537] = 8'h00;
Memory[17536] = 8'hB8;
Memory[17543] = 8'h00;
Memory[17542] = 8'h00;
Memory[17541] = 8'h00;
Memory[17540] = 8'h92;
Memory[17547] = 8'h00;
Memory[17546] = 8'h00;
Memory[17545] = 8'h00;
Memory[17544] = 8'hA4;
Memory[17551] = 8'h00;
Memory[17550] = 8'h00;
Memory[17549] = 8'h01;
Memory[17548] = 8'h15;
Memory[17555] = 8'h00;
Memory[17554] = 8'h00;
Memory[17553] = 8'h01;
Memory[17552] = 8'h25;
Memory[17559] = 8'h00;
Memory[17558] = 8'h00;
Memory[17557] = 8'h01;
Memory[17556] = 8'h71;
Memory[17563] = 8'h00;
Memory[17562] = 8'h00;
Memory[17561] = 8'h01;
Memory[17560] = 8'hB8;
Memory[17567] = 8'h00;
Memory[17566] = 8'h00;
Memory[17565] = 8'h00;
Memory[17564] = 8'hDC;
Memory[17571] = 8'h00;
Memory[17570] = 8'h00;
Memory[17569] = 8'h00;
Memory[17568] = 8'hF6;
Memory[17575] = 8'h00;
Memory[17574] = 8'h00;
Memory[17573] = 8'h00;
Memory[17572] = 8'hC3;
Memory[17579] = 8'h00;
Memory[17578] = 8'h00;
Memory[17577] = 8'h00;
Memory[17576] = 8'hDC;
Memory[17583] = 8'h00;
Memory[17582] = 8'h00;
Memory[17581] = 8'h00;
Memory[17580] = 8'hB8;
Memory[17587] = 8'h00;
Memory[17586] = 8'h00;
Memory[17585] = 8'h00;
Memory[17584] = 8'h92;
Memory[17591] = 8'h00;
Memory[17590] = 8'h00;
Memory[17589] = 8'h01;
Memory[17588] = 8'h25;
Memory[17595] = 8'h00;
Memory[17594] = 8'h00;
Memory[17593] = 8'h01;
Memory[17592] = 8'h15;
Memory[17599] = 8'h00;
Memory[17598] = 8'h00;
Memory[17597] = 8'h01;
Memory[17596] = 8'h25;
Memory[17603] = 8'h00;
Memory[17602] = 8'h00;
Memory[17601] = 8'h01;
Memory[17600] = 8'h15;
Memory[17607] = 8'h00;
Memory[17606] = 8'h00;
Memory[17605] = 8'h01;
Memory[17604] = 8'h25;
Memory[17611] = 8'h00;
Memory[17610] = 8'h00;
Memory[17609] = 8'h00;
Memory[17608] = 8'h92;
Memory[17615] = 8'h00;
Memory[17614] = 8'h00;
Memory[17613] = 8'h00;
Memory[17612] = 8'h8A;
Memory[17619] = 8'h00;
Memory[17618] = 8'h00;
Memory[17617] = 8'h00;
Memory[17616] = 8'hDC;
Memory[17623] = 8'h00;
Memory[17622] = 8'h00;
Memory[17621] = 8'h00;
Memory[17620] = 8'hA4;
Memory[17627] = 8'h00;
Memory[17626] = 8'h00;
Memory[17625] = 8'h00;
Memory[17624] = 8'hB8;
Memory[17631] = 8'h00;
Memory[17630] = 8'h00;
Memory[17629] = 8'h00;
Memory[17628] = 8'h92;
Memory[17635] = 8'h00;
Memory[17634] = 8'h00;
Memory[17633] = 8'h01;
Memory[17632] = 8'h25;
Memory[17639] = 8'h00;
Memory[17638] = 8'h00;
Memory[17637] = 8'h01;
Memory[17636] = 8'h15;
Memory[17643] = 8'h00;
Memory[17642] = 8'h00;
Memory[17641] = 8'h00;
Memory[17640] = 8'hF6;
Memory[17647] = 8'h00;
Memory[17646] = 8'h00;
Memory[17645] = 8'h01;
Memory[17644] = 8'h15;
Memory[17651] = 8'h00;
Memory[17650] = 8'h00;
Memory[17649] = 8'h01;
Memory[17648] = 8'h71;
Memory[17655] = 8'h00;
Memory[17654] = 8'h00;
Memory[17653] = 8'h01;
Memory[17652] = 8'hB8;
Memory[17659] = 8'h00;
Memory[17658] = 8'h00;
Memory[17657] = 8'h01;
Memory[17656] = 8'hED;
Memory[17663] = 8'h00;
Memory[17662] = 8'h00;
Memory[17661] = 8'h01;
Memory[17660] = 8'h87;
Memory[17667] = 8'h00;
Memory[17666] = 8'h00;
Memory[17665] = 8'h01;
Memory[17664] = 8'h71;
Memory[17671] = 8'h00;
Memory[17670] = 8'h00;
Memory[17669] = 8'h01;
Memory[17668] = 8'h49;
Memory[17675] = 8'h00;
Memory[17674] = 8'h00;
Memory[17673] = 8'h01;
Memory[17672] = 8'h87;
Memory[17679] = 8'h00;
Memory[17678] = 8'h00;
Memory[17677] = 8'h01;
Memory[17676] = 8'h71;
Memory[17683] = 8'h00;
Memory[17682] = 8'h00;
Memory[17681] = 8'h01;
Memory[17680] = 8'h49;
Memory[17687] = 8'h00;
Memory[17686] = 8'h00;
Memory[17685] = 8'h01;
Memory[17684] = 8'h25;
Memory[17691] = 8'h00;
Memory[17690] = 8'h00;
Memory[17689] = 8'h01;
Memory[17688] = 8'h15;
Memory[17695] = 8'h00;
Memory[17694] = 8'h00;
Memory[17693] = 8'h00;
Memory[17692] = 8'hF6;
Memory[17699] = 8'h00;
Memory[17698] = 8'h00;
Memory[17697] = 8'h00;
Memory[17696] = 8'hDC;
Memory[17703] = 8'h00;
Memory[17702] = 8'h00;
Memory[17701] = 8'h00;
Memory[17700] = 8'hC3;
Memory[17707] = 8'h00;
Memory[17706] = 8'h00;
Memory[17705] = 8'h00;
Memory[17704] = 8'hB8;
Memory[17711] = 8'h00;
Memory[17710] = 8'h00;
Memory[17709] = 8'h00;
Memory[17708] = 8'hA4;
Memory[17715] = 8'h00;
Memory[17714] = 8'h00;
Memory[17713] = 8'h00;
Memory[17712] = 8'hC3;
Memory[17719] = 8'h00;
Memory[17718] = 8'h00;
Memory[17717] = 8'h00;
Memory[17716] = 8'hB8;
Memory[17723] = 8'h00;
Memory[17722] = 8'h00;
Memory[17721] = 8'h00;
Memory[17720] = 8'hA4;
Memory[17727] = 8'h00;
Memory[17726] = 8'h00;
Memory[17725] = 8'h00;
Memory[17724] = 8'h92;
Memory[17731] = 8'h00;
Memory[17730] = 8'h00;
Memory[17729] = 8'h00;
Memory[17728] = 8'hA4;
Memory[17735] = 8'h00;
Memory[17734] = 8'h00;
Memory[17733] = 8'h00;
Memory[17732] = 8'hB8;
Memory[17739] = 8'h00;
Memory[17738] = 8'h00;
Memory[17737] = 8'h00;
Memory[17736] = 8'hC3;
Memory[17743] = 8'h00;
Memory[17742] = 8'h00;
Memory[17741] = 8'h00;
Memory[17740] = 8'hDC;
Memory[17747] = 8'h00;
Memory[17746] = 8'h00;
Memory[17745] = 8'h00;
Memory[17744] = 8'hA4;
Memory[17751] = 8'h00;
Memory[17750] = 8'h00;
Memory[17749] = 8'h00;
Memory[17748] = 8'hDC;
Memory[17755] = 8'h00;
Memory[17754] = 8'h00;
Memory[17753] = 8'h00;
Memory[17752] = 8'hC3;
Memory[17759] = 8'h00;
Memory[17758] = 8'h00;
Memory[17757] = 8'h00;
Memory[17756] = 8'hB8;
Memory[17763] = 8'h00;
Memory[17762] = 8'h00;
Memory[17761] = 8'h00;
Memory[17760] = 8'hF6;
Memory[17767] = 8'h00;
Memory[17766] = 8'h00;
Memory[17765] = 8'h00;
Memory[17764] = 8'hDC;
Memory[17771] = 8'h00;
Memory[17770] = 8'h00;
Memory[17769] = 8'h00;
Memory[17768] = 8'hC3;
Memory[17775] = 8'h00;
Memory[17774] = 8'h00;
Memory[17773] = 8'h00;
Memory[17772] = 8'hDC;
Memory[17779] = 8'h00;
Memory[17778] = 8'h00;
Memory[17777] = 8'h00;
Memory[17776] = 8'hC3;
Memory[17783] = 8'h00;
Memory[17782] = 8'h00;
Memory[17781] = 8'h00;
Memory[17780] = 8'hB8;
Memory[17787] = 8'h00;
Memory[17786] = 8'h00;
Memory[17785] = 8'h00;
Memory[17784] = 8'hA4;
Memory[17791] = 8'h00;
Memory[17790] = 8'h00;
Memory[17789] = 8'h00;
Memory[17788] = 8'h92;
Memory[17795] = 8'h00;
Memory[17794] = 8'h00;
Memory[17793] = 8'h00;
Memory[17792] = 8'hF6;
Memory[17799] = 8'h00;
Memory[17798] = 8'h00;
Memory[17797] = 8'h01;
Memory[17796] = 8'h15;
Memory[17803] = 8'h00;
Memory[17802] = 8'h00;
Memory[17801] = 8'h01;
Memory[17800] = 8'h25;
Memory[17807] = 8'h00;
Memory[17806] = 8'h00;
Memory[17805] = 8'h01;
Memory[17804] = 8'h15;
Memory[17811] = 8'h00;
Memory[17810] = 8'h00;
Memory[17809] = 8'h00;
Memory[17808] = 8'hF6;
Memory[17815] = 8'h00;
Memory[17814] = 8'h00;
Memory[17813] = 8'h00;
Memory[17812] = 8'hDC;
Memory[17819] = 8'h00;
Memory[17818] = 8'h00;
Memory[17817] = 8'h00;
Memory[17816] = 8'hC3;
Memory[17823] = 8'h00;
Memory[17822] = 8'h00;
Memory[17821] = 8'h00;
Memory[17820] = 8'hB8;
Memory[17827] = 8'h00;
Memory[17826] = 8'h00;
Memory[17825] = 8'h00;
Memory[17824] = 8'hA4;
Memory[17831] = 8'h00;
Memory[17830] = 8'h00;
Memory[17829] = 8'h00;
Memory[17828] = 8'hF6;
Memory[17835] = 8'h00;
Memory[17834] = 8'h00;
Memory[17833] = 8'h00;
Memory[17832] = 8'hDC;
Memory[17839] = 8'h00;
Memory[17838] = 8'h00;
Memory[17837] = 8'h00;
Memory[17836] = 8'hF6;
Memory[17843] = 8'h00;
Memory[17842] = 8'h00;
Memory[17841] = 8'h00;
Memory[17840] = 8'hDC;
Memory[17847] = 8'h00;
Memory[17846] = 8'h00;
Memory[17845] = 8'h00;
Memory[17844] = 8'hC3;
Memory[17851] = 8'h00;
Memory[17850] = 8'h00;
Memory[17849] = 8'h00;
Memory[17848] = 8'hB8;
Memory[17855] = 8'h00;
Memory[17854] = 8'h00;
Memory[17853] = 8'h01;
Memory[17852] = 8'h71;
Memory[17859] = 8'h00;
Memory[17858] = 8'h00;
Memory[17857] = 8'h01;
Memory[17856] = 8'h49;
Memory[17863] = 8'h00;
Memory[17862] = 8'h00;
Memory[17861] = 8'h00;
Memory[17860] = 8'h00;
Memory[17867] = 8'h00;
Memory[17866] = 8'h00;
Memory[17865] = 8'h01;
Memory[17864] = 8'h25;
Memory[17871] = 8'h00;
Memory[17870] = 8'h00;
Memory[17869] = 8'h01;
Memory[17868] = 8'h71;
Memory[17875] = 8'h00;
Memory[17874] = 8'h00;
Memory[17873] = 8'h01;
Memory[17872] = 8'hED;
Memory[17879] = 8'h00;
Memory[17878] = 8'h00;
Memory[17877] = 8'h01;
Memory[17876] = 8'hB8;
Memory[17883] = 8'h00;
Memory[17882] = 8'h00;
Memory[17881] = 8'h01;
Memory[17880] = 8'hED;
Memory[17887] = 8'h00;
Memory[17886] = 8'h00;
Memory[17885] = 8'h02;
Memory[17884] = 8'h2A;
Memory[17891] = 8'h00;
Memory[17890] = 8'h00;
Memory[17889] = 8'h02;
Memory[17888] = 8'h4B;
Memory[17895] = 8'h00;
Memory[17894] = 8'h00;
Memory[17893] = 8'h01;
Memory[17892] = 8'h25;
Memory[17899] = 8'h00;
Memory[17898] = 8'h00;
Memory[17897] = 8'h01;
Memory[17896] = 8'h15;
Memory[17903] = 8'h00;
Memory[17902] = 8'h00;
Memory[17901] = 8'h00;
Memory[17900] = 8'h00;
Memory[17907] = 8'h00;
Memory[17906] = 8'h00;
Memory[17905] = 8'h00;
Memory[17904] = 8'hF6;
Memory[17911] = 8'h00;
Memory[17910] = 8'h00;
Memory[17909] = 8'h01;
Memory[17908] = 8'h25;
Memory[17915] = 8'h00;
Memory[17914] = 8'h00;
Memory[17913] = 8'h01;
Memory[17912] = 8'h87;
Memory[17919] = 8'h00;
Memory[17918] = 8'h00;
Memory[17917] = 8'h01;
Memory[17916] = 8'h49;
Memory[17923] = 8'h00;
Memory[17922] = 8'h00;
Memory[17921] = 8'h01;
Memory[17920] = 8'hB8;
Memory[17927] = 8'h00;
Memory[17926] = 8'h00;
Memory[17925] = 8'h01;
Memory[17924] = 8'h71;
Memory[17931] = 8'h00;
Memory[17930] = 8'h00;
Memory[17929] = 8'h01;
Memory[17928] = 8'h87;
Memory[17935] = 8'h00;
Memory[17934] = 8'h00;
Memory[17933] = 8'h01;
Memory[17932] = 8'hB8;
Memory[17939] = 8'h00;
Memory[17938] = 8'h00;
Memory[17937] = 8'h01;
Memory[17936] = 8'h71;
Memory[17943] = 8'h00;
Memory[17942] = 8'h00;
Memory[17941] = 8'h01;
Memory[17940] = 8'h87;
Memory[17947] = 8'h00;
Memory[17946] = 8'h00;
Memory[17945] = 8'h01;
Memory[17944] = 8'hB8;
Memory[17951] = 8'h00;
Memory[17950] = 8'h00;
Memory[17949] = 8'h00;
Memory[17948] = 8'hDC;
Memory[17955] = 8'h00;
Memory[17954] = 8'h00;
Memory[17953] = 8'h00;
Memory[17952] = 8'hF6;
Memory[17959] = 8'h00;
Memory[17958] = 8'h00;
Memory[17957] = 8'h01;
Memory[17956] = 8'h15;
Memory[17963] = 8'h00;
Memory[17962] = 8'h00;
Memory[17961] = 8'h01;
Memory[17960] = 8'h25;
Memory[17967] = 8'h00;
Memory[17966] = 8'h00;
Memory[17965] = 8'h01;
Memory[17964] = 8'h49;
Memory[17971] = 8'h00;
Memory[17970] = 8'h00;
Memory[17969] = 8'h01;
Memory[17968] = 8'h71;
Memory[17975] = 8'h00;
Memory[17974] = 8'h00;
Memory[17973] = 8'h01;
Memory[17972] = 8'h87;
Memory[17979] = 8'h00;
Memory[17978] = 8'h00;
Memory[17977] = 8'h01;
Memory[17976] = 8'h71;
Memory[17983] = 8'h00;
Memory[17982] = 8'h00;
Memory[17981] = 8'h01;
Memory[17980] = 8'h25;
Memory[17987] = 8'h00;
Memory[17986] = 8'h00;
Memory[17985] = 8'h01;
Memory[17984] = 8'h49;
Memory[17991] = 8'h00;
Memory[17990] = 8'h00;
Memory[17989] = 8'h01;
Memory[17988] = 8'h71;
Memory[17995] = 8'h00;
Memory[17994] = 8'h00;
Memory[17993] = 8'h00;
Memory[17992] = 8'hB8;
Memory[17999] = 8'h00;
Memory[17998] = 8'h00;
Memory[17997] = 8'h00;
Memory[17996] = 8'hC3;
Memory[18003] = 8'h00;
Memory[18002] = 8'h00;
Memory[18001] = 8'h00;
Memory[18000] = 8'hDC;
Memory[18007] = 8'h00;
Memory[18006] = 8'h00;
Memory[18005] = 8'h00;
Memory[18004] = 8'hF6;
Memory[18011] = 8'h00;
Memory[18010] = 8'h00;
Memory[18009] = 8'h00;
Memory[18008] = 8'hDC;
Memory[18015] = 8'h00;
Memory[18014] = 8'h00;
Memory[18013] = 8'h00;
Memory[18012] = 8'hC3;
Memory[18019] = 8'h00;
Memory[18018] = 8'h00;
Memory[18017] = 8'h00;
Memory[18016] = 8'hDC;
Memory[18023] = 8'h00;
Memory[18022] = 8'h00;
Memory[18021] = 8'h00;
Memory[18020] = 8'hB8;
Memory[18027] = 8'h00;
Memory[18026] = 8'h00;
Memory[18025] = 8'h00;
Memory[18024] = 8'hC3;
Memory[18031] = 8'h00;
Memory[18030] = 8'h00;
Memory[18029] = 8'h00;
Memory[18028] = 8'hDC;
Memory[18035] = 8'h00;
Memory[18034] = 8'h00;
Memory[18033] = 8'h00;
Memory[18032] = 8'hC3;
Memory[18039] = 8'h00;
Memory[18038] = 8'h00;
Memory[18037] = 8'h00;
Memory[18036] = 8'hF6;
Memory[18043] = 8'h00;
Memory[18042] = 8'h00;
Memory[18041] = 8'h00;
Memory[18040] = 8'hDC;
Memory[18047] = 8'h00;
Memory[18046] = 8'h00;
Memory[18045] = 8'h00;
Memory[18044] = 8'hC3;
Memory[18051] = 8'h00;
Memory[18050] = 8'h00;
Memory[18049] = 8'h00;
Memory[18048] = 8'hB8;
Memory[18055] = 8'h00;
Memory[18054] = 8'h00;
Memory[18053] = 8'h00;
Memory[18052] = 8'hA4;
Memory[18059] = 8'h00;
Memory[18058] = 8'h00;
Memory[18057] = 8'h00;
Memory[18056] = 8'hB8;
Memory[18063] = 8'h00;
Memory[18062] = 8'h00;
Memory[18061] = 8'h00;
Memory[18060] = 8'hA4;
Memory[18067] = 8'h00;
Memory[18066] = 8'h00;
Memory[18065] = 8'h00;
Memory[18064] = 8'h92;
Memory[18071] = 8'h00;
Memory[18070] = 8'h00;
Memory[18069] = 8'h00;
Memory[18068] = 8'hA4;
Memory[18075] = 8'h00;
Memory[18074] = 8'h00;
Memory[18073] = 8'h00;
Memory[18072] = 8'hB8;
Memory[18079] = 8'h00;
Memory[18078] = 8'h00;
Memory[18077] = 8'h00;
Memory[18076] = 8'hC3;
Memory[18083] = 8'h00;
Memory[18082] = 8'h00;
Memory[18081] = 8'h00;
Memory[18080] = 8'hDC;
Memory[18087] = 8'h00;
Memory[18086] = 8'h00;
Memory[18085] = 8'h00;
Memory[18084] = 8'hF6;
Memory[18091] = 8'h00;
Memory[18090] = 8'h00;
Memory[18089] = 8'h00;
Memory[18088] = 8'hC3;
Memory[18095] = 8'h00;
Memory[18094] = 8'h00;
Memory[18093] = 8'h00;
Memory[18092] = 8'hF6;
Memory[18099] = 8'h00;
Memory[18098] = 8'h00;
Memory[18097] = 8'h00;
Memory[18096] = 8'hDC;
Memory[18103] = 8'h00;
Memory[18102] = 8'h00;
Memory[18101] = 8'h00;
Memory[18100] = 8'hF6;
Memory[18107] = 8'h00;
Memory[18106] = 8'h00;
Memory[18105] = 8'h01;
Memory[18104] = 8'h15;
Memory[18111] = 8'h00;
Memory[18110] = 8'h00;
Memory[18109] = 8'h01;
Memory[18108] = 8'h25;
Memory[18115] = 8'h00;
Memory[18114] = 8'h00;
Memory[18113] = 8'h00;
Memory[18112] = 8'hDC;
Memory[18119] = 8'h00;
Memory[18118] = 8'h00;
Memory[18117] = 8'h00;
Memory[18116] = 8'hF6;
Memory[18123] = 8'h00;
Memory[18122] = 8'h00;
Memory[18121] = 8'h01;
Memory[18120] = 8'h15;
Memory[18127] = 8'h00;
Memory[18126] = 8'h00;
Memory[18125] = 8'h01;
Memory[18124] = 8'h25;
Memory[18131] = 8'h00;
Memory[18130] = 8'h00;
Memory[18129] = 8'h01;
Memory[18128] = 8'h49;
Memory[18135] = 8'h00;
Memory[18134] = 8'h00;
Memory[18133] = 8'h01;
Memory[18132] = 8'h71;
Memory[18139] = 8'h00;
Memory[18138] = 8'h00;
Memory[18137] = 8'h01;
Memory[18136] = 8'h87;
Memory[18143] = 8'h00;
Memory[18142] = 8'h00;
Memory[18141] = 8'h01;
Memory[18140] = 8'hB8;
Memory[18147] = 8'h00;
Memory[18146] = 8'h00;
Memory[18145] = 8'h01;
Memory[18144] = 8'h71;
Memory[18151] = 8'h00;
Memory[18150] = 8'h00;
Memory[18149] = 8'h01;
Memory[18148] = 8'h25;
Memory[18155] = 8'h00;
Memory[18154] = 8'h00;
Memory[18153] = 8'h01;
Memory[18152] = 8'h49;
Memory[18159] = 8'h00;
Memory[18158] = 8'h00;
Memory[18157] = 8'h01;
Memory[18156] = 8'h71;
Memory[18163] = 8'h00;
Memory[18162] = 8'h00;
Memory[18161] = 8'h01;
Memory[18160] = 8'h49;
Memory[18167] = 8'h00;
Memory[18166] = 8'h00;
Memory[18165] = 8'h01;
Memory[18164] = 8'h25;
Memory[18171] = 8'h00;
Memory[18170] = 8'h00;
Memory[18169] = 8'h01;
Memory[18168] = 8'h49;
Memory[18175] = 8'h00;
Memory[18174] = 8'h00;
Memory[18173] = 8'h00;
Memory[18172] = 8'hDC;
Memory[18179] = 8'h00;
Memory[18178] = 8'h00;
Memory[18177] = 8'h00;
Memory[18176] = 8'hF6;
Memory[18183] = 8'h00;
Memory[18182] = 8'h00;
Memory[18181] = 8'h01;
Memory[18180] = 8'h49;
Memory[18187] = 8'h00;
Memory[18186] = 8'h00;
Memory[18185] = 8'h01;
Memory[18184] = 8'h71;
Memory[18191] = 8'h00;
Memory[18190] = 8'h00;
Memory[18189] = 8'h01;
Memory[18188] = 8'h49;
Memory[18195] = 8'h00;
Memory[18194] = 8'h00;
Memory[18193] = 8'h01;
Memory[18192] = 8'h25;
Memory[18199] = 8'h00;
Memory[18198] = 8'h00;
Memory[18197] = 8'h01;
Memory[18196] = 8'h15;
Memory[18203] = 8'h00;
Memory[18202] = 8'h00;
Memory[18201] = 8'h01;
Memory[18200] = 8'h25;
Memory[18207] = 8'h00;
Memory[18206] = 8'h00;
Memory[18205] = 8'h00;
Memory[18204] = 8'hF6;
Memory[18211] = 8'h00;
Memory[18210] = 8'h00;
Memory[18209] = 8'h01;
Memory[18208] = 8'h15;
Memory[18215] = 8'h00;
Memory[18214] = 8'h00;
Memory[18213] = 8'h01;
Memory[18212] = 8'h25;
Memory[18219] = 8'h00;
Memory[18218] = 8'h00;
Memory[18217] = 8'h00;
Memory[18216] = 8'h92;
Memory[18223] = 8'h00;
Memory[18222] = 8'h00;
Memory[18221] = 8'h00;
Memory[18220] = 8'hA4;
Memory[18227] = 8'h00;
Memory[18226] = 8'h00;
Memory[18225] = 8'h00;
Memory[18224] = 8'hB8;
Memory[18231] = 8'h00;
Memory[18230] = 8'h00;
Memory[18229] = 8'h00;
Memory[18228] = 8'hC3;
Memory[18235] = 8'h00;
Memory[18234] = 8'h00;
Memory[18233] = 8'h00;
Memory[18232] = 8'hB8;
Memory[18239] = 8'h00;
Memory[18238] = 8'h00;
Memory[18237] = 8'h00;
Memory[18236] = 8'hA4;
Memory[18243] = 8'h00;
Memory[18242] = 8'h00;
Memory[18241] = 8'h00;
Memory[18240] = 8'hB8;
Memory[18247] = 8'h00;
Memory[18246] = 8'h00;
Memory[18245] = 8'h01;
Memory[18244] = 8'h25;
Memory[18251] = 8'h00;
Memory[18250] = 8'h00;
Memory[18249] = 8'h01;
Memory[18248] = 8'h15;
Memory[18255] = 8'h00;
Memory[18254] = 8'h00;
Memory[18253] = 8'h01;
Memory[18252] = 8'h25;
Memory[18259] = 8'h00;
Memory[18258] = 8'h00;
Memory[18257] = 8'h00;
Memory[18256] = 8'hF6;
Memory[18263] = 8'h00;
Memory[18262] = 8'h00;
Memory[18261] = 8'h01;
Memory[18260] = 8'h25;
Memory[18267] = 8'h00;
Memory[18266] = 8'h00;
Memory[18265] = 8'h01;
Memory[18264] = 8'h15;
Memory[18271] = 8'h00;
Memory[18270] = 8'h00;
Memory[18269] = 8'h00;
Memory[18268] = 8'hF6;
Memory[18275] = 8'h00;
Memory[18274] = 8'h00;
Memory[18273] = 8'h00;
Memory[18272] = 8'hDC;
Memory[18279] = 8'h00;
Memory[18278] = 8'h00;
Memory[18277] = 8'h00;
Memory[18276] = 8'hC3;
Memory[18283] = 8'h00;
Memory[18282] = 8'h00;
Memory[18281] = 8'h00;
Memory[18280] = 8'hDC;
Memory[18287] = 8'h00;
Memory[18286] = 8'h00;
Memory[18285] = 8'h00;
Memory[18284] = 8'hC3;
Memory[18291] = 8'h00;
Memory[18290] = 8'h00;
Memory[18289] = 8'h00;
Memory[18288] = 8'hB8;
Memory[18295] = 8'h00;
Memory[18294] = 8'h00;
Memory[18293] = 8'h00;
Memory[18292] = 8'hC3;
Memory[18299] = 8'h00;
Memory[18298] = 8'h00;
Memory[18297] = 8'h00;
Memory[18296] = 8'hDC;
Memory[18303] = 8'h00;
Memory[18302] = 8'h00;
Memory[18301] = 8'h00;
Memory[18300] = 8'hF6;
Memory[18307] = 8'h00;
Memory[18306] = 8'h00;
Memory[18305] = 8'h01;
Memory[18304] = 8'h15;
Memory[18311] = 8'h00;
Memory[18310] = 8'h00;
Memory[18309] = 8'h01;
Memory[18308] = 8'h25;
Memory[18315] = 8'h00;
Memory[18314] = 8'h00;
Memory[18313] = 8'h00;
Memory[18312] = 8'hF6;
Memory[18319] = 8'h00;
Memory[18318] = 8'h00;
Memory[18317] = 8'h01;
Memory[18316] = 8'h25;
Memory[18323] = 8'h00;
Memory[18322] = 8'h00;
Memory[18321] = 8'h01;
Memory[18320] = 8'h15;
Memory[18327] = 8'h00;
Memory[18326] = 8'h00;
Memory[18325] = 8'h01;
Memory[18324] = 8'h25;
Memory[18331] = 8'h00;
Memory[18330] = 8'h00;
Memory[18329] = 8'h01;
Memory[18328] = 8'h15;
Memory[18335] = 8'h00;
Memory[18334] = 8'h00;
Memory[18333] = 8'h00;
Memory[18332] = 8'hF6;
Memory[18339] = 8'h00;
Memory[18338] = 8'h00;
Memory[18337] = 8'h01;
Memory[18336] = 8'h15;
Memory[18343] = 8'h00;
Memory[18342] = 8'h00;
Memory[18341] = 8'h01;
Memory[18340] = 8'h25;
Memory[18347] = 8'h00;
Memory[18346] = 8'h00;
Memory[18345] = 8'h01;
Memory[18344] = 8'h49;
Memory[18351] = 8'h00;
Memory[18350] = 8'h00;
Memory[18349] = 8'h01;
Memory[18348] = 8'h25;
Memory[18355] = 8'h00;
Memory[18354] = 8'h00;
Memory[18353] = 8'h01;
Memory[18352] = 8'h15;
Memory[18359] = 8'h00;
Memory[18358] = 8'h00;
Memory[18357] = 8'h01;
Memory[18356] = 8'h25;
Memory[18363] = 8'h00;
Memory[18362] = 8'h00;
Memory[18361] = 8'h00;
Memory[18360] = 8'hF6;
Memory[18367] = 8'h00;
Memory[18366] = 8'h00;
Memory[18365] = 8'h01;
Memory[18364] = 8'h15;
Memory[18371] = 8'h00;
Memory[18370] = 8'h00;
Memory[18369] = 8'h01;
Memory[18368] = 8'hB8;
Memory[18375] = 8'h00;
Memory[18374] = 8'h00;
Memory[18373] = 8'h01;
Memory[18372] = 8'h71;
Memory[18379] = 8'h00;
Memory[18378] = 8'h00;
Memory[18377] = 8'h01;
Memory[18376] = 8'h87;
Memory[18383] = 8'h00;
Memory[18382] = 8'h00;
Memory[18381] = 8'h01;
Memory[18380] = 8'hB8;
Memory[18387] = 8'h00;
Memory[18386] = 8'h00;
Memory[18385] = 8'h01;
Memory[18384] = 8'h71;
Memory[18391] = 8'h00;
Memory[18390] = 8'h00;
Memory[18389] = 8'h01;
Memory[18388] = 8'h87;
Memory[18395] = 8'h00;
Memory[18394] = 8'h00;
Memory[18393] = 8'h01;
Memory[18392] = 8'hB8;
Memory[18399] = 8'h00;
Memory[18398] = 8'h00;
Memory[18397] = 8'h00;
Memory[18396] = 8'hDC;
Memory[18403] = 8'h00;
Memory[18402] = 8'h00;
Memory[18401] = 8'h00;
Memory[18400] = 8'hF6;
Memory[18407] = 8'h00;
Memory[18406] = 8'h00;
Memory[18405] = 8'h01;
Memory[18404] = 8'h15;
Memory[18411] = 8'h00;
Memory[18410] = 8'h00;
Memory[18409] = 8'h01;
Memory[18408] = 8'h25;
Memory[18415] = 8'h00;
Memory[18414] = 8'h00;
Memory[18413] = 8'h01;
Memory[18412] = 8'h49;
Memory[18419] = 8'h00;
Memory[18418] = 8'h00;
Memory[18417] = 8'h01;
Memory[18416] = 8'h71;
Memory[18423] = 8'h00;
Memory[18422] = 8'h00;
Memory[18421] = 8'h01;
Memory[18420] = 8'h87;
Memory[18427] = 8'h00;
Memory[18426] = 8'h00;
Memory[18425] = 8'h01;
Memory[18424] = 8'h71;
Memory[18431] = 8'h00;
Memory[18430] = 8'h00;
Memory[18429] = 8'h01;
Memory[18428] = 8'h25;
Memory[18435] = 8'h00;
Memory[18434] = 8'h00;
Memory[18433] = 8'h01;
Memory[18432] = 8'h49;
Memory[18439] = 8'h00;
Memory[18438] = 8'h00;
Memory[18437] = 8'h01;
Memory[18436] = 8'h71;
Memory[18443] = 8'h00;
Memory[18442] = 8'h00;
Memory[18441] = 8'h00;
Memory[18440] = 8'hB8;
Memory[18447] = 8'h00;
Memory[18446] = 8'h00;
Memory[18445] = 8'h00;
Memory[18444] = 8'hC3;
Memory[18451] = 8'h00;
Memory[18450] = 8'h00;
Memory[18449] = 8'h00;
Memory[18448] = 8'hDC;
Memory[18455] = 8'h00;
Memory[18454] = 8'h00;
Memory[18453] = 8'h00;
Memory[18452] = 8'hF6;
Memory[18459] = 8'h00;
Memory[18458] = 8'h00;
Memory[18457] = 8'h00;
Memory[18456] = 8'hDC;
Memory[18463] = 8'h00;
Memory[18462] = 8'h00;
Memory[18461] = 8'h00;
Memory[18460] = 8'hC3;
Memory[18467] = 8'h00;
Memory[18466] = 8'h00;
Memory[18465] = 8'h00;
Memory[18464] = 8'hDC;
Memory[18471] = 8'h00;
Memory[18470] = 8'h00;
Memory[18469] = 8'h00;
Memory[18468] = 8'hB8;
Memory[18475] = 8'h00;
Memory[18474] = 8'h00;
Memory[18473] = 8'h00;
Memory[18472] = 8'hC3;
Memory[18479] = 8'h00;
Memory[18478] = 8'h00;
Memory[18477] = 8'h00;
Memory[18476] = 8'hDC;
Memory[18483] = 8'h00;
Memory[18482] = 8'h00;
Memory[18481] = 8'h00;
Memory[18480] = 8'hC3;
Memory[18487] = 8'h00;
Memory[18486] = 8'h00;
Memory[18485] = 8'h00;
Memory[18484] = 8'hF6;
Memory[18491] = 8'h00;
Memory[18490] = 8'h00;
Memory[18489] = 8'h00;
Memory[18488] = 8'hDC;
Memory[18495] = 8'h00;
Memory[18494] = 8'h00;
Memory[18493] = 8'h00;
Memory[18492] = 8'hC3;
Memory[18499] = 8'h00;
Memory[18498] = 8'h00;
Memory[18497] = 8'h00;
Memory[18496] = 8'hB8;
Memory[18503] = 8'h00;
Memory[18502] = 8'h00;
Memory[18501] = 8'h00;
Memory[18500] = 8'hA4;
Memory[18507] = 8'h00;
Memory[18506] = 8'h00;
Memory[18505] = 8'h00;
Memory[18504] = 8'hB8;
Memory[18511] = 8'h00;
Memory[18510] = 8'h00;
Memory[18509] = 8'h00;
Memory[18508] = 8'hA4;
Memory[18515] = 8'h00;
Memory[18514] = 8'h00;
Memory[18513] = 8'h00;
Memory[18512] = 8'h92;
Memory[18519] = 8'h00;
Memory[18518] = 8'h00;
Memory[18517] = 8'h00;
Memory[18516] = 8'hA4;
Memory[18523] = 8'h00;
Memory[18522] = 8'h00;
Memory[18521] = 8'h00;
Memory[18520] = 8'hB8;
Memory[18527] = 8'h00;
Memory[18526] = 8'h00;
Memory[18525] = 8'h00;
Memory[18524] = 8'hC3;
Memory[18531] = 8'h00;
Memory[18530] = 8'h00;
Memory[18529] = 8'h00;
Memory[18528] = 8'hDC;
Memory[18535] = 8'h00;
Memory[18534] = 8'h00;
Memory[18533] = 8'h00;
Memory[18532] = 8'hF6;
Memory[18539] = 8'h00;
Memory[18538] = 8'h00;
Memory[18537] = 8'h00;
Memory[18536] = 8'hC3;
Memory[18543] = 8'h00;
Memory[18542] = 8'h00;
Memory[18541] = 8'h00;
Memory[18540] = 8'hF6;
Memory[18547] = 8'h00;
Memory[18546] = 8'h00;
Memory[18545] = 8'h00;
Memory[18544] = 8'hDC;
Memory[18551] = 8'h00;
Memory[18550] = 8'h00;
Memory[18549] = 8'h00;
Memory[18548] = 8'hF6;
Memory[18555] = 8'h00;
Memory[18554] = 8'h00;
Memory[18553] = 8'h01;
Memory[18552] = 8'h15;
Memory[18559] = 8'h00;
Memory[18558] = 8'h00;
Memory[18557] = 8'h01;
Memory[18556] = 8'h25;
Memory[18563] = 8'h00;
Memory[18562] = 8'h00;
Memory[18561] = 8'h00;
Memory[18560] = 8'hDC;
Memory[18567] = 8'h00;
Memory[18566] = 8'h00;
Memory[18565] = 8'h00;
Memory[18564] = 8'hF6;
Memory[18571] = 8'h00;
Memory[18570] = 8'h00;
Memory[18569] = 8'h01;
Memory[18568] = 8'h15;
Memory[18575] = 8'h00;
Memory[18574] = 8'h00;
Memory[18573] = 8'h01;
Memory[18572] = 8'h25;
Memory[18579] = 8'h00;
Memory[18578] = 8'h00;
Memory[18577] = 8'h01;
Memory[18576] = 8'h49;
Memory[18583] = 8'h00;
Memory[18582] = 8'h00;
Memory[18581] = 8'h01;
Memory[18580] = 8'h71;
Memory[18587] = 8'h00;
Memory[18586] = 8'h00;
Memory[18585] = 8'h01;
Memory[18584] = 8'h87;
Memory[18591] = 8'h00;
Memory[18590] = 8'h00;
Memory[18589] = 8'h01;
Memory[18588] = 8'hB8;
Memory[18595] = 8'h00;
Memory[18594] = 8'h00;
Memory[18593] = 8'h01;
Memory[18592] = 8'h71;
Memory[18599] = 8'h00;
Memory[18598] = 8'h00;
Memory[18597] = 8'h01;
Memory[18596] = 8'h25;
Memory[18603] = 8'h00;
Memory[18602] = 8'h00;
Memory[18601] = 8'h01;
Memory[18600] = 8'h49;
Memory[18607] = 8'h00;
Memory[18606] = 8'h00;
Memory[18605] = 8'h01;
Memory[18604] = 8'h71;
Memory[18611] = 8'h00;
Memory[18610] = 8'h00;
Memory[18609] = 8'h01;
Memory[18608] = 8'h49;
Memory[18615] = 8'h00;
Memory[18614] = 8'h00;
Memory[18613] = 8'h01;
Memory[18612] = 8'h25;
Memory[18619] = 8'h00;
Memory[18618] = 8'h00;
Memory[18617] = 8'h01;
Memory[18616] = 8'h49;
Memory[18623] = 8'h00;
Memory[18622] = 8'h00;
Memory[18621] = 8'h00;
Memory[18620] = 8'hDC;
Memory[18627] = 8'h00;
Memory[18626] = 8'h00;
Memory[18625] = 8'h00;
Memory[18624] = 8'hF6;
Memory[18631] = 8'h00;
Memory[18630] = 8'h00;
Memory[18629] = 8'h01;
Memory[18628] = 8'h49;
Memory[18635] = 8'h00;
Memory[18634] = 8'h00;
Memory[18633] = 8'h01;
Memory[18632] = 8'h71;
Memory[18639] = 8'h00;
Memory[18638] = 8'h00;
Memory[18637] = 8'h01;
Memory[18636] = 8'h49;
Memory[18643] = 8'h00;
Memory[18642] = 8'h00;
Memory[18641] = 8'h01;
Memory[18640] = 8'h25;
Memory[18647] = 8'h00;
Memory[18646] = 8'h00;
Memory[18645] = 8'h01;
Memory[18644] = 8'h15;
Memory[18651] = 8'h00;
Memory[18650] = 8'h00;
Memory[18649] = 8'h01;
Memory[18648] = 8'h25;
Memory[18655] = 8'h00;
Memory[18654] = 8'h00;
Memory[18653] = 8'h00;
Memory[18652] = 8'hF6;
Memory[18659] = 8'h00;
Memory[18658] = 8'h00;
Memory[18657] = 8'h01;
Memory[18656] = 8'h15;
Memory[18663] = 8'h00;
Memory[18662] = 8'h00;
Memory[18661] = 8'h01;
Memory[18660] = 8'h25;
Memory[18667] = 8'h00;
Memory[18666] = 8'h00;
Memory[18665] = 8'h00;
Memory[18664] = 8'h92;
Memory[18671] = 8'h00;
Memory[18670] = 8'h00;
Memory[18669] = 8'h00;
Memory[18668] = 8'hA4;
Memory[18675] = 8'h00;
Memory[18674] = 8'h00;
Memory[18673] = 8'h00;
Memory[18672] = 8'hB8;
Memory[18679] = 8'h00;
Memory[18678] = 8'h00;
Memory[18677] = 8'h00;
Memory[18676] = 8'hC3;
Memory[18683] = 8'h00;
Memory[18682] = 8'h00;
Memory[18681] = 8'h00;
Memory[18680] = 8'hB8;
Memory[18687] = 8'h00;
Memory[18686] = 8'h00;
Memory[18685] = 8'h00;
Memory[18684] = 8'hA4;
Memory[18691] = 8'h00;
Memory[18690] = 8'h00;
Memory[18689] = 8'h00;
Memory[18688] = 8'hB8;
Memory[18695] = 8'h00;
Memory[18694] = 8'h00;
Memory[18693] = 8'h01;
Memory[18692] = 8'h25;
Memory[18699] = 8'h00;
Memory[18698] = 8'h00;
Memory[18697] = 8'h01;
Memory[18696] = 8'h15;
Memory[18703] = 8'h00;
Memory[18702] = 8'h00;
Memory[18701] = 8'h01;
Memory[18700] = 8'h25;
Memory[18707] = 8'h00;
Memory[18706] = 8'h00;
Memory[18705] = 8'h00;
Memory[18704] = 8'hF6;
Memory[18711] = 8'h00;
Memory[18710] = 8'h00;
Memory[18709] = 8'h01;
Memory[18708] = 8'h25;
Memory[18715] = 8'h00;
Memory[18714] = 8'h00;
Memory[18713] = 8'h01;
Memory[18712] = 8'h15;
Memory[18719] = 8'h00;
Memory[18718] = 8'h00;
Memory[18717] = 8'h00;
Memory[18716] = 8'hF6;
Memory[18723] = 8'h00;
Memory[18722] = 8'h00;
Memory[18721] = 8'h00;
Memory[18720] = 8'hDC;
Memory[18727] = 8'h00;
Memory[18726] = 8'h00;
Memory[18725] = 8'h00;
Memory[18724] = 8'hC3;
Memory[18731] = 8'h00;
Memory[18730] = 8'h00;
Memory[18729] = 8'h00;
Memory[18728] = 8'hDC;
Memory[18735] = 8'h00;
Memory[18734] = 8'h00;
Memory[18733] = 8'h00;
Memory[18732] = 8'hC3;
Memory[18739] = 8'h00;
Memory[18738] = 8'h00;
Memory[18737] = 8'h00;
Memory[18736] = 8'hB8;
Memory[18743] = 8'h00;
Memory[18742] = 8'h00;
Memory[18741] = 8'h00;
Memory[18740] = 8'hC3;
Memory[18747] = 8'h00;
Memory[18746] = 8'h00;
Memory[18745] = 8'h00;
Memory[18744] = 8'hDC;
Memory[18751] = 8'h00;
Memory[18750] = 8'h00;
Memory[18749] = 8'h00;
Memory[18748] = 8'hF6;
Memory[18755] = 8'h00;
Memory[18754] = 8'h00;
Memory[18753] = 8'h01;
Memory[18752] = 8'h15;
Memory[18759] = 8'h00;
Memory[18758] = 8'h00;
Memory[18757] = 8'h01;
Memory[18756] = 8'h25;
Memory[18763] = 8'h00;
Memory[18762] = 8'h00;
Memory[18761] = 8'h00;
Memory[18760] = 8'hF6;
Memory[18767] = 8'h00;
Memory[18766] = 8'h00;
Memory[18765] = 8'h01;
Memory[18764] = 8'h25;
Memory[18771] = 8'h00;
Memory[18770] = 8'h00;
Memory[18769] = 8'h01;
Memory[18768] = 8'h15;
Memory[18775] = 8'h00;
Memory[18774] = 8'h00;
Memory[18773] = 8'h01;
Memory[18772] = 8'h25;
Memory[18779] = 8'h00;
Memory[18778] = 8'h00;
Memory[18777] = 8'h01;
Memory[18776] = 8'h15;
Memory[18783] = 8'h00;
Memory[18782] = 8'h00;
Memory[18781] = 8'h00;
Memory[18780] = 8'hF6;
Memory[18787] = 8'h00;
Memory[18786] = 8'h00;
Memory[18785] = 8'h01;
Memory[18784] = 8'h15;
Memory[18791] = 8'h00;
Memory[18790] = 8'h00;
Memory[18789] = 8'h01;
Memory[18788] = 8'h25;
Memory[18795] = 8'h00;
Memory[18794] = 8'h00;
Memory[18793] = 8'h01;
Memory[18792] = 8'h49;
Memory[18799] = 8'h00;
Memory[18798] = 8'h00;
Memory[18797] = 8'h01;
Memory[18796] = 8'h25;
Memory[18803] = 8'h00;
Memory[18802] = 8'h00;
Memory[18801] = 8'h01;
Memory[18800] = 8'h15;
Memory[18807] = 8'h00;
Memory[18806] = 8'h00;
Memory[18805] = 8'h01;
Memory[18804] = 8'h25;
Memory[18811] = 8'h00;
Memory[18810] = 8'h00;
Memory[18809] = 8'h00;
Memory[18808] = 8'hF6;
Memory[18815] = 8'h00;
Memory[18814] = 8'h00;
Memory[18813] = 8'h01;
Memory[18812] = 8'h15;
Memory[18819] = 8'h00;
Memory[18818] = 8'h00;
Memory[18817] = 8'h00;
Memory[18816] = 8'hB8;
Memory[18823] = 8'h00;
Memory[18822] = 8'h00;
Memory[18821] = 8'h01;
Memory[18820] = 8'h71;
Memory[18827] = 8'h00;
Memory[18826] = 8'h00;
Memory[18825] = 8'h01;
Memory[18824] = 8'h87;
Memory[18831] = 8'h00;
Memory[18830] = 8'h00;
Memory[18829] = 8'h01;
Memory[18828] = 8'h71;
Memory[18835] = 8'h00;
Memory[18834] = 8'h00;
Memory[18833] = 8'h01;
Memory[18832] = 8'h49;
Memory[18839] = 8'h00;
Memory[18838] = 8'h00;
Memory[18837] = 8'h01;
Memory[18836] = 8'h25;
Memory[18843] = 8'h00;
Memory[18842] = 8'h00;
Memory[18841] = 8'h01;
Memory[18840] = 8'h49;
Memory[18847] = 8'h00;
Memory[18846] = 8'h00;
Memory[18845] = 8'h01;
Memory[18844] = 8'h25;
Memory[18851] = 8'h00;
Memory[18850] = 8'h00;
Memory[18849] = 8'h01;
Memory[18848] = 8'h15;
Memory[18855] = 8'h00;
Memory[18854] = 8'h00;
Memory[18853] = 8'h00;
Memory[18852] = 8'hF6;
Memory[18859] = 8'h00;
Memory[18858] = 8'h00;
Memory[18857] = 8'h01;
Memory[18856] = 8'h25;
Memory[18863] = 8'h00;
Memory[18862] = 8'h00;
Memory[18861] = 8'h01;
Memory[18860] = 8'h15;
Memory[18867] = 8'h00;
Memory[18866] = 8'h00;
Memory[18865] = 8'h00;
Memory[18864] = 8'hF6;
Memory[18871] = 8'h00;
Memory[18870] = 8'h00;
Memory[18869] = 8'h01;
Memory[18868] = 8'h15;
Memory[18875] = 8'h00;
Memory[18874] = 8'h00;
Memory[18873] = 8'h00;
Memory[18872] = 8'hDC;
Memory[18879] = 8'h00;
Memory[18878] = 8'h00;
Memory[18877] = 8'h01;
Memory[18876] = 8'hB8;
Memory[18883] = 8'h00;
Memory[18882] = 8'h00;
Memory[18881] = 8'h01;
Memory[18880] = 8'hED;
Memory[18887] = 8'h00;
Memory[18886] = 8'h00;
Memory[18885] = 8'h01;
Memory[18884] = 8'hB8;
Memory[18891] = 8'h00;
Memory[18890] = 8'h00;
Memory[18889] = 8'h01;
Memory[18888] = 8'h87;
Memory[18895] = 8'h00;
Memory[18894] = 8'h00;
Memory[18893] = 8'h01;
Memory[18892] = 8'h71;
Memory[18899] = 8'h00;
Memory[18898] = 8'h00;
Memory[18897] = 8'h01;
Memory[18896] = 8'h87;
Memory[18903] = 8'h00;
Memory[18902] = 8'h00;
Memory[18901] = 8'h01;
Memory[18900] = 8'h71;
Memory[18907] = 8'h00;
Memory[18906] = 8'h00;
Memory[18905] = 8'h01;
Memory[18904] = 8'h49;
Memory[18911] = 8'h00;
Memory[18910] = 8'h00;
Memory[18909] = 8'h01;
Memory[18908] = 8'h25;
Memory[18915] = 8'h00;
Memory[18914] = 8'h00;
Memory[18913] = 8'h01;
Memory[18912] = 8'h15;
Memory[18919] = 8'h00;
Memory[18918] = 8'h00;
Memory[18917] = 8'h00;
Memory[18916] = 8'hF6;
Memory[18923] = 8'h00;
Memory[18922] = 8'h00;
Memory[18921] = 8'h01;
Memory[18920] = 8'h15;
Memory[18927] = 8'h00;
Memory[18926] = 8'h00;
Memory[18925] = 8'h00;
Memory[18924] = 8'hDC;
Memory[18931] = 8'h00;
Memory[18930] = 8'h00;
Memory[18929] = 8'h00;
Memory[18928] = 8'hC3;
Memory[18935] = 8'h00;
Memory[18934] = 8'h00;
Memory[18933] = 8'h01;
Memory[18932] = 8'h25;
Memory[18939] = 8'h00;
Memory[18938] = 8'h00;
Memory[18937] = 8'h01;
Memory[18936] = 8'h15;
Memory[18943] = 8'h00;
Memory[18942] = 8'h00;
Memory[18941] = 8'h00;
Memory[18940] = 8'hB8;
Memory[18947] = 8'h00;
Memory[18946] = 8'h00;
Memory[18945] = 8'h01;
Memory[18944] = 8'h71;
Memory[18951] = 8'h00;
Memory[18950] = 8'h00;
Memory[18949] = 8'h01;
Memory[18948] = 8'h87;
Memory[18955] = 8'h00;
Memory[18954] = 8'h00;
Memory[18953] = 8'h01;
Memory[18952] = 8'h71;
Memory[18959] = 8'h00;
Memory[18958] = 8'h00;
Memory[18957] = 8'h01;
Memory[18956] = 8'h49;
Memory[18963] = 8'h00;
Memory[18962] = 8'h00;
Memory[18961] = 8'h01;
Memory[18960] = 8'h25;
Memory[18967] = 8'h00;
Memory[18966] = 8'h00;
Memory[18965] = 8'h01;
Memory[18964] = 8'h49;
Memory[18971] = 8'h00;
Memory[18970] = 8'h00;
Memory[18969] = 8'h01;
Memory[18968] = 8'h25;
Memory[18975] = 8'h00;
Memory[18974] = 8'h00;
Memory[18973] = 8'h01;
Memory[18972] = 8'h15;
Memory[18979] = 8'h00;
Memory[18978] = 8'h00;
Memory[18977] = 8'h00;
Memory[18976] = 8'hF6;
Memory[18983] = 8'h00;
Memory[18982] = 8'h00;
Memory[18981] = 8'h01;
Memory[18980] = 8'h25;
Memory[18987] = 8'h00;
Memory[18986] = 8'h00;
Memory[18985] = 8'h01;
Memory[18984] = 8'h15;
Memory[18991] = 8'h00;
Memory[18990] = 8'h00;
Memory[18989] = 8'h00;
Memory[18988] = 8'hF6;
Memory[18995] = 8'h00;
Memory[18994] = 8'h00;
Memory[18993] = 8'h01;
Memory[18992] = 8'h15;
Memory[18999] = 8'h00;
Memory[18998] = 8'h00;
Memory[18997] = 8'h00;
Memory[18996] = 8'hDC;
Memory[19003] = 8'h00;
Memory[19002] = 8'h00;
Memory[19001] = 8'h01;
Memory[19000] = 8'hB8;
Memory[19007] = 8'h00;
Memory[19006] = 8'h00;
Memory[19005] = 8'h01;
Memory[19004] = 8'hED;
Memory[19011] = 8'h00;
Memory[19010] = 8'h00;
Memory[19009] = 8'h01;
Memory[19008] = 8'hB8;
Memory[19015] = 8'h00;
Memory[19014] = 8'h00;
Memory[19013] = 8'h01;
Memory[19012] = 8'h87;
Memory[19019] = 8'h00;
Memory[19018] = 8'h00;
Memory[19017] = 8'h01;
Memory[19016] = 8'h71;
Memory[19023] = 8'h00;
Memory[19022] = 8'h00;
Memory[19021] = 8'h01;
Memory[19020] = 8'h87;
Memory[19027] = 8'h00;
Memory[19026] = 8'h00;
Memory[19025] = 8'h01;
Memory[19024] = 8'h71;
Memory[19031] = 8'h00;
Memory[19030] = 8'h00;
Memory[19029] = 8'h01;
Memory[19028] = 8'h49;
Memory[19035] = 8'h00;
Memory[19034] = 8'h00;
Memory[19033] = 8'h01;
Memory[19032] = 8'h25;
Memory[19039] = 8'h00;
Memory[19038] = 8'h00;
Memory[19037] = 8'h01;
Memory[19036] = 8'h15;
Memory[19043] = 8'h00;
Memory[19042] = 8'h00;
Memory[19041] = 8'h00;
Memory[19040] = 8'hF6;
Memory[19047] = 8'h00;
Memory[19046] = 8'h00;
Memory[19045] = 8'h01;
Memory[19044] = 8'h15;
Memory[19051] = 8'h00;
Memory[19050] = 8'h00;
Memory[19049] = 8'h00;
Memory[19048] = 8'hDC;
Memory[19055] = 8'h00;
Memory[19054] = 8'h00;
Memory[19053] = 8'h00;
Memory[19052] = 8'hC3;
Memory[19059] = 8'h00;
Memory[19058] = 8'h00;
Memory[19057] = 8'h01;
Memory[19056] = 8'h25;
Memory[19063] = 8'h00;
Memory[19062] = 8'h00;
Memory[19061] = 8'h01;
Memory[19060] = 8'h15;
Memory[19067] = 8'h00;
Memory[19066] = 8'h00;
Memory[19065] = 8'h01;
Memory[19064] = 8'h71;
Memory[19071] = 8'h00;
Memory[19070] = 8'h00;
Memory[19069] = 8'h01;
Memory[19068] = 8'h49;
Memory[19075] = 8'h00;
Memory[19074] = 8'h00;
Memory[19073] = 8'h01;
Memory[19072] = 8'h25;
Memory[19079] = 8'h00;
Memory[19078] = 8'h00;
Memory[19077] = 8'h01;
Memory[19076] = 8'h15;
Memory[19083] = 8'h00;
Memory[19082] = 8'h00;
Memory[19081] = 8'h00;
Memory[19080] = 8'hF6;
Memory[19087] = 8'h00;
Memory[19086] = 8'h00;
Memory[19085] = 8'h00;
Memory[19084] = 8'hDC;
Memory[19091] = 8'h00;
Memory[19090] = 8'h00;
Memory[19089] = 8'h00;
Memory[19088] = 8'hF6;
Memory[19095] = 8'h00;
Memory[19094] = 8'h00;
Memory[19093] = 8'h01;
Memory[19092] = 8'h15;
Memory[19099] = 8'h00;
Memory[19098] = 8'h00;
Memory[19097] = 8'h01;
Memory[19096] = 8'h25;
Memory[19103] = 8'h00;
Memory[19102] = 8'h00;
Memory[19101] = 8'h01;
Memory[19100] = 8'h15;
Memory[19107] = 8'h00;
Memory[19106] = 8'h00;
Memory[19105] = 8'h00;
Memory[19104] = 8'hF6;
Memory[19111] = 8'h00;
Memory[19110] = 8'h00;
Memory[19109] = 8'h00;
Memory[19108] = 8'hDC;
Memory[19115] = 8'h00;
Memory[19114] = 8'h00;
Memory[19113] = 8'h00;
Memory[19112] = 8'hF6;
Memory[19119] = 8'h00;
Memory[19118] = 8'h00;
Memory[19117] = 8'h01;
Memory[19116] = 8'h25;
Memory[19123] = 8'h00;
Memory[19122] = 8'h00;
Memory[19121] = 8'h01;
Memory[19120] = 8'h71;
Memory[19127] = 8'h00;
Memory[19126] = 8'h00;
Memory[19125] = 8'h01;
Memory[19124] = 8'h25;
Memory[19131] = 8'h00;
Memory[19130] = 8'h00;
Memory[19129] = 8'h00;
Memory[19128] = 8'hF6;
Memory[19135] = 8'h00;
Memory[19134] = 8'h00;
Memory[19133] = 8'h01;
Memory[19132] = 8'h15;
Memory[19139] = 8'h00;
Memory[19138] = 8'h00;
Memory[19137] = 8'h01;
Memory[19136] = 8'h25;
Memory[19143] = 8'h00;
Memory[19142] = 8'h00;
Memory[19141] = 8'h00;
Memory[19140] = 8'h00;
Memory[19147] = 8'h00;
Memory[19146] = 8'h0D;
Memory[19145] = 8'h21;
Memory[19144] = 8'h83;
Memory[19151] = 8'h00;
Memory[19150] = 8'h3B;
Memory[19149] = 8'h2A;
Memory[19148] = 8'h23;
Memory[19155] = 8'h12;
Memory[19154] = 8'h40;
Memory[19153] = 8'h20;
Memory[19152] = 8'h6F;
Memory[19159] = 8'h00;
Memory[19158] = 8'h4D;
Memory[19157] = 8'h21;
Memory[19156] = 8'h83;
Memory[19163] = 8'h00;
Memory[19162] = 8'h3B;
Memory[19161] = 8'h2A;
Memory[19160] = 8'h23;
Memory[19167] = 8'h12;
Memory[19166] = 8'h40;
Memory[19165] = 8'h20;
Memory[19164] = 8'h6F;
Memory[19171] = 8'h00;
Memory[19170] = 8'h8D;
Memory[19169] = 8'h21;
Memory[19168] = 8'h83;
Memory[19175] = 8'h00;
Memory[19174] = 8'h3B;
Memory[19173] = 8'h2A;
Memory[19172] = 8'h23;
Memory[19179] = 8'h12;
Memory[19178] = 8'h40;
Memory[19177] = 8'h20;
Memory[19176] = 8'h6F;
Memory[19183] = 8'h00;
Memory[19182] = 8'hCD;
Memory[19181] = 8'h21;
Memory[19180] = 8'h83;
Memory[19187] = 8'h00;
Memory[19186] = 8'h3B;
Memory[19185] = 8'h2A;
Memory[19184] = 8'h23;
Memory[19191] = 8'h12;
Memory[19190] = 8'h40;
Memory[19189] = 8'h20;
Memory[19188] = 8'h6F;
Memory[19195] = 8'h01;
Memory[19194] = 8'h0D;
Memory[19193] = 8'h21;
Memory[19192] = 8'h83;
Memory[19199] = 8'h00;
Memory[19198] = 8'h3B;
Memory[19197] = 8'h2A;
Memory[19196] = 8'h23;
Memory[19203] = 8'h12;
Memory[19202] = 8'h40;
Memory[19201] = 8'h20;
Memory[19200] = 8'h6F;
Memory[19207] = 8'h01;
Memory[19206] = 8'h4D;
Memory[19205] = 8'h21;
Memory[19204] = 8'h83;
Memory[19211] = 8'h00;
Memory[19210] = 8'h3B;
Memory[19209] = 8'h2A;
Memory[19208] = 8'h23;
Memory[19215] = 8'h12;
Memory[19214] = 8'h40;
Memory[19213] = 8'h20;
Memory[19212] = 8'h6F;
Memory[19219] = 8'h01;
Memory[19218] = 8'h8D;
Memory[19217] = 8'h21;
Memory[19216] = 8'h83;
Memory[19223] = 8'h00;
Memory[19222] = 8'h3B;
Memory[19221] = 8'h2A;
Memory[19220] = 8'h23;
Memory[19227] = 8'h12;
Memory[19226] = 8'h40;
Memory[19225] = 8'h20;
Memory[19224] = 8'h6F;
Memory[19231] = 8'h01;
Memory[19230] = 8'hCD;
Memory[19229] = 8'h21;
Memory[19228] = 8'h83;
Memory[19235] = 8'h00;
Memory[19234] = 8'h3B;
Memory[19233] = 8'h2A;
Memory[19232] = 8'h23;
Memory[19239] = 8'h12;
Memory[19238] = 8'h40;
Memory[19237] = 8'h20;
Memory[19236] = 8'h6F;
Memory[19243] = 8'h02;
Memory[19242] = 8'h0D;
Memory[19241] = 8'h21;
Memory[19240] = 8'h83;
Memory[19247] = 8'h00;
Memory[19246] = 8'h3B;
Memory[19245] = 8'h2A;
Memory[19244] = 8'h23;
Memory[19251] = 8'h12;
Memory[19250] = 8'h40;
Memory[19249] = 8'h20;
Memory[19248] = 8'h6F;
Memory[19255] = 8'h02;
Memory[19254] = 8'h4D;
Memory[19253] = 8'h21;
Memory[19252] = 8'h83;
Memory[19259] = 8'h00;
Memory[19258] = 8'h3B;
Memory[19257] = 8'h2A;
Memory[19256] = 8'h23;
Memory[19263] = 8'h12;
Memory[19262] = 8'h40;
Memory[19261] = 8'h20;
Memory[19260] = 8'h6F;
Memory[19267] = 8'h02;
Memory[19266] = 8'h8D;
Memory[19265] = 8'h21;
Memory[19264] = 8'h83;
Memory[19271] = 8'h00;
Memory[19270] = 8'h3B;
Memory[19269] = 8'h2A;
Memory[19268] = 8'h23;
Memory[19275] = 8'h12;
Memory[19274] = 8'h40;
Memory[19273] = 8'h20;
Memory[19272] = 8'h6F;
Memory[19279] = 8'h02;
Memory[19278] = 8'hCD;
Memory[19277] = 8'h21;
Memory[19276] = 8'h83;
Memory[19283] = 8'h00;
Memory[19282] = 8'h3B;
Memory[19281] = 8'h2A;
Memory[19280] = 8'h23;
Memory[19287] = 8'h12;
Memory[19286] = 8'h40;
Memory[19285] = 8'h20;
Memory[19284] = 8'h6F;
Memory[19291] = 8'h03;
Memory[19290] = 8'h0D;
Memory[19289] = 8'h21;
Memory[19288] = 8'h83;
Memory[19295] = 8'h00;
Memory[19294] = 8'h3B;
Memory[19293] = 8'h2A;
Memory[19292] = 8'h23;
Memory[19299] = 8'h12;
Memory[19298] = 8'h40;
Memory[19297] = 8'h20;
Memory[19296] = 8'h6F;
Memory[19303] = 8'h03;
Memory[19302] = 8'h4D;
Memory[19301] = 8'h21;
Memory[19300] = 8'h83;
Memory[19307] = 8'h00;
Memory[19306] = 8'h3B;
Memory[19305] = 8'h2A;
Memory[19304] = 8'h23;
Memory[19311] = 8'h12;
Memory[19310] = 8'h40;
Memory[19309] = 8'h20;
Memory[19308] = 8'h6F;
Memory[19315] = 8'h03;
Memory[19314] = 8'h8D;
Memory[19313] = 8'h21;
Memory[19312] = 8'h83;
Memory[19319] = 8'h00;
Memory[19318] = 8'h3B;
Memory[19317] = 8'h2A;
Memory[19316] = 8'h23;
Memory[19323] = 8'h12;
Memory[19322] = 8'h40;
Memory[19321] = 8'h20;
Memory[19320] = 8'h6F;
Memory[19327] = 8'h03;
Memory[19326] = 8'hCD;
Memory[19325] = 8'h21;
Memory[19324] = 8'h83;
Memory[19331] = 8'h00;
Memory[19330] = 8'h3B;
Memory[19329] = 8'h2A;
Memory[19328] = 8'h23;
Memory[19335] = 8'h12;
Memory[19334] = 8'h40;
Memory[19333] = 8'h20;
Memory[19332] = 8'h6F;
Memory[19339] = 8'h04;
Memory[19338] = 8'h0D;
Memory[19337] = 8'h21;
Memory[19336] = 8'h83;
Memory[19343] = 8'h00;
Memory[19342] = 8'h3B;
Memory[19341] = 8'h2A;
Memory[19340] = 8'h23;
Memory[19347] = 8'h12;
Memory[19346] = 8'h40;
Memory[19345] = 8'h20;
Memory[19344] = 8'h6F;
Memory[19351] = 8'h04;
Memory[19350] = 8'h4D;
Memory[19349] = 8'h21;
Memory[19348] = 8'h83;
Memory[19355] = 8'h00;
Memory[19354] = 8'h3B;
Memory[19353] = 8'h2A;
Memory[19352] = 8'h23;
Memory[19359] = 8'h12;
Memory[19358] = 8'h40;
Memory[19357] = 8'h20;
Memory[19356] = 8'h6F;
Memory[19363] = 8'h04;
Memory[19362] = 8'h8D;
Memory[19361] = 8'h21;
Memory[19360] = 8'h83;
Memory[19367] = 8'h00;
Memory[19366] = 8'h3B;
Memory[19365] = 8'h2A;
Memory[19364] = 8'h23;
Memory[19371] = 8'h12;
Memory[19370] = 8'h40;
Memory[19369] = 8'h20;
Memory[19368] = 8'h6F;
Memory[19375] = 8'h04;
Memory[19374] = 8'hCD;
Memory[19373] = 8'h21;
Memory[19372] = 8'h83;
Memory[19379] = 8'h00;
Memory[19378] = 8'h3B;
Memory[19377] = 8'h2A;
Memory[19376] = 8'h23;
Memory[19383] = 8'h12;
Memory[19382] = 8'h40;
Memory[19381] = 8'h20;
Memory[19380] = 8'h6F;
Memory[19387] = 8'h05;
Memory[19386] = 8'h0D;
Memory[19385] = 8'h21;
Memory[19384] = 8'h83;
Memory[19391] = 8'h00;
Memory[19390] = 8'h3B;
Memory[19389] = 8'h2A;
Memory[19388] = 8'h23;
Memory[19395] = 8'h12;
Memory[19394] = 8'h40;
Memory[19393] = 8'h20;
Memory[19392] = 8'h6F;
Memory[19399] = 8'h05;
Memory[19398] = 8'h4D;
Memory[19397] = 8'h21;
Memory[19396] = 8'h83;
Memory[19403] = 8'h00;
Memory[19402] = 8'h3B;
Memory[19401] = 8'h2A;
Memory[19400] = 8'h23;
Memory[19407] = 8'h12;
Memory[19406] = 8'h40;
Memory[19405] = 8'h20;
Memory[19404] = 8'h6F;
Memory[19411] = 8'h05;
Memory[19410] = 8'h8D;
Memory[19409] = 8'h21;
Memory[19408] = 8'h83;
Memory[19415] = 8'h00;
Memory[19414] = 8'h3B;
Memory[19413] = 8'h2A;
Memory[19412] = 8'h23;
Memory[19419] = 8'h12;
Memory[19418] = 8'h40;
Memory[19417] = 8'h20;
Memory[19416] = 8'h6F;
Memory[19423] = 8'h05;
Memory[19422] = 8'hCD;
Memory[19421] = 8'h21;
Memory[19420] = 8'h83;
Memory[19427] = 8'h00;
Memory[19426] = 8'h3B;
Memory[19425] = 8'h2A;
Memory[19424] = 8'h23;
Memory[19431] = 8'h12;
Memory[19430] = 8'h40;
Memory[19429] = 8'h20;
Memory[19428] = 8'h6F;
Memory[19435] = 8'h06;
Memory[19434] = 8'h0D;
Memory[19433] = 8'h21;
Memory[19432] = 8'h83;
Memory[19439] = 8'h00;
Memory[19438] = 8'h3B;
Memory[19437] = 8'h2A;
Memory[19436] = 8'h23;
Memory[19443] = 8'h12;
Memory[19442] = 8'h40;
Memory[19441] = 8'h20;
Memory[19440] = 8'h6F;
Memory[19447] = 8'h06;
Memory[19446] = 8'h4D;
Memory[19445] = 8'h21;
Memory[19444] = 8'h83;
Memory[19451] = 8'h00;
Memory[19450] = 8'h3B;
Memory[19449] = 8'h2A;
Memory[19448] = 8'h23;
Memory[19455] = 8'h12;
Memory[19454] = 8'h40;
Memory[19453] = 8'h20;
Memory[19452] = 8'h6F;
Memory[19459] = 8'h06;
Memory[19458] = 8'h8D;
Memory[19457] = 8'h21;
Memory[19456] = 8'h83;
Memory[19463] = 8'h00;
Memory[19462] = 8'h3B;
Memory[19461] = 8'h2A;
Memory[19460] = 8'h23;
Memory[19467] = 8'h12;
Memory[19466] = 8'h40;
Memory[19465] = 8'h20;
Memory[19464] = 8'h6F;
Memory[19471] = 8'h06;
Memory[19470] = 8'hCD;
Memory[19469] = 8'h21;
Memory[19468] = 8'h83;
Memory[19475] = 8'h00;
Memory[19474] = 8'h3B;
Memory[19473] = 8'h2A;
Memory[19472] = 8'h23;
Memory[19479] = 8'h12;
Memory[19478] = 8'h40;
Memory[19477] = 8'h20;
Memory[19476] = 8'h6F;
Memory[19483] = 8'h07;
Memory[19482] = 8'h0D;
Memory[19481] = 8'h21;
Memory[19480] = 8'h83;
Memory[19487] = 8'h00;
Memory[19486] = 8'h3B;
Memory[19485] = 8'h2A;
Memory[19484] = 8'h23;
Memory[19491] = 8'h12;
Memory[19490] = 8'h40;
Memory[19489] = 8'h20;
Memory[19488] = 8'h6F;
Memory[19495] = 8'h07;
Memory[19494] = 8'h4D;
Memory[19493] = 8'h21;
Memory[19492] = 8'h83;
Memory[19499] = 8'h00;
Memory[19498] = 8'h3B;
Memory[19497] = 8'h2A;
Memory[19496] = 8'h23;
Memory[19503] = 8'h12;
Memory[19502] = 8'h40;
Memory[19501] = 8'h20;
Memory[19500] = 8'h6F;
Memory[19507] = 8'h07;
Memory[19506] = 8'h8D;
Memory[19505] = 8'h21;
Memory[19504] = 8'h83;
Memory[19511] = 8'h00;
Memory[19510] = 8'h3B;
Memory[19509] = 8'h2A;
Memory[19508] = 8'h23;
Memory[19515] = 8'h12;
Memory[19514] = 8'h40;
Memory[19513] = 8'h20;
Memory[19512] = 8'h6F;
Memory[19519] = 8'h07;
Memory[19518] = 8'hCD;
Memory[19517] = 8'h21;
Memory[19516] = 8'h83;
Memory[19523] = 8'h00;
Memory[19522] = 8'h3B;
Memory[19521] = 8'h2A;
Memory[19520] = 8'h23;
Memory[19527] = 8'h12;
Memory[19526] = 8'h40;
Memory[19525] = 8'h20;
Memory[19524] = 8'h6F;
Memory[19531] = 8'h08;
Memory[19530] = 8'h0D;
Memory[19529] = 8'h21;
Memory[19528] = 8'h83;
Memory[19535] = 8'h00;
Memory[19534] = 8'h3B;
Memory[19533] = 8'h2A;
Memory[19532] = 8'h23;
Memory[19539] = 8'h12;
Memory[19538] = 8'h40;
Memory[19537] = 8'h20;
Memory[19536] = 8'h6F;
Memory[19543] = 8'h08;
Memory[19542] = 8'h4D;
Memory[19541] = 8'h21;
Memory[19540] = 8'h83;
Memory[19547] = 8'h00;
Memory[19546] = 8'h3B;
Memory[19545] = 8'h2A;
Memory[19544] = 8'h23;
Memory[19551] = 8'h12;
Memory[19550] = 8'h40;
Memory[19549] = 8'h20;
Memory[19548] = 8'h6F;
Memory[19555] = 8'h08;
Memory[19554] = 8'h8D;
Memory[19553] = 8'h21;
Memory[19552] = 8'h83;
Memory[19559] = 8'h00;
Memory[19558] = 8'h3B;
Memory[19557] = 8'h2A;
Memory[19556] = 8'h23;
Memory[19563] = 8'h12;
Memory[19562] = 8'h40;
Memory[19561] = 8'h20;
Memory[19560] = 8'h6F;
Memory[19567] = 8'h08;
Memory[19566] = 8'hCD;
Memory[19565] = 8'h21;
Memory[19564] = 8'h83;
Memory[19571] = 8'h00;
Memory[19570] = 8'h3B;
Memory[19569] = 8'h2A;
Memory[19568] = 8'h23;
Memory[19575] = 8'h12;
Memory[19574] = 8'h40;
Memory[19573] = 8'h20;
Memory[19572] = 8'h6F;
Memory[19579] = 8'h09;
Memory[19578] = 8'h0D;
Memory[19577] = 8'h21;
Memory[19576] = 8'h83;
Memory[19583] = 8'h00;
Memory[19582] = 8'h3B;
Memory[19581] = 8'h2A;
Memory[19580] = 8'h23;
Memory[19587] = 8'h12;
Memory[19586] = 8'h40;
Memory[19585] = 8'h20;
Memory[19584] = 8'h6F;
Memory[19591] = 8'h09;
Memory[19590] = 8'h4D;
Memory[19589] = 8'h21;
Memory[19588] = 8'h83;
Memory[19595] = 8'h00;
Memory[19594] = 8'h3B;
Memory[19593] = 8'h2A;
Memory[19592] = 8'h23;
Memory[19599] = 8'h12;
Memory[19598] = 8'h40;
Memory[19597] = 8'h20;
Memory[19596] = 8'h6F;
Memory[19603] = 8'h09;
Memory[19602] = 8'h8D;
Memory[19601] = 8'h21;
Memory[19600] = 8'h83;
Memory[19607] = 8'h00;
Memory[19606] = 8'h3B;
Memory[19605] = 8'h2A;
Memory[19604] = 8'h23;
Memory[19611] = 8'h12;
Memory[19610] = 8'h40;
Memory[19609] = 8'h20;
Memory[19608] = 8'h6F;
Memory[19615] = 8'h09;
Memory[19614] = 8'hCD;
Memory[19613] = 8'h21;
Memory[19612] = 8'h83;
Memory[19619] = 8'h00;
Memory[19618] = 8'h3B;
Memory[19617] = 8'h2A;
Memory[19616] = 8'h23;
Memory[19623] = 8'h12;
Memory[19622] = 8'h40;
Memory[19621] = 8'h20;
Memory[19620] = 8'h6F;
Memory[19627] = 8'h0A;
Memory[19626] = 8'h0D;
Memory[19625] = 8'h21;
Memory[19624] = 8'h83;
Memory[19631] = 8'h00;
Memory[19630] = 8'h3B;
Memory[19629] = 8'h2A;
Memory[19628] = 8'h23;
Memory[19635] = 8'h12;
Memory[19634] = 8'h40;
Memory[19633] = 8'h20;
Memory[19632] = 8'h6F;
Memory[19639] = 8'h0A;
Memory[19638] = 8'h4D;
Memory[19637] = 8'h21;
Memory[19636] = 8'h83;
Memory[19643] = 8'h00;
Memory[19642] = 8'h3B;
Memory[19641] = 8'h2A;
Memory[19640] = 8'h23;
Memory[19647] = 8'h12;
Memory[19646] = 8'h40;
Memory[19645] = 8'h20;
Memory[19644] = 8'h6F;
Memory[19651] = 8'h0A;
Memory[19650] = 8'h8D;
Memory[19649] = 8'h21;
Memory[19648] = 8'h83;
Memory[19655] = 8'h00;
Memory[19654] = 8'h3B;
Memory[19653] = 8'h2A;
Memory[19652] = 8'h23;
Memory[19659] = 8'h12;
Memory[19658] = 8'h40;
Memory[19657] = 8'h20;
Memory[19656] = 8'h6F;
Memory[19663] = 8'h0A;
Memory[19662] = 8'hCD;
Memory[19661] = 8'h21;
Memory[19660] = 8'h83;
Memory[19667] = 8'h00;
Memory[19666] = 8'h3B;
Memory[19665] = 8'h2A;
Memory[19664] = 8'h23;
Memory[19671] = 8'h12;
Memory[19670] = 8'h40;
Memory[19669] = 8'h20;
Memory[19668] = 8'h6F;
Memory[19675] = 8'h0B;
Memory[19674] = 8'h0D;
Memory[19673] = 8'h21;
Memory[19672] = 8'h83;
Memory[19679] = 8'h00;
Memory[19678] = 8'h3B;
Memory[19677] = 8'h2A;
Memory[19676] = 8'h23;
Memory[19683] = 8'h12;
Memory[19682] = 8'h40;
Memory[19681] = 8'h20;
Memory[19680] = 8'h6F;
Memory[19687] = 8'h0B;
Memory[19686] = 8'h4D;
Memory[19685] = 8'h21;
Memory[19684] = 8'h83;
Memory[19691] = 8'h00;
Memory[19690] = 8'h3B;
Memory[19689] = 8'h2A;
Memory[19688] = 8'h23;
Memory[19695] = 8'h12;
Memory[19694] = 8'h40;
Memory[19693] = 8'h20;
Memory[19692] = 8'h6F;
Memory[19699] = 8'h0B;
Memory[19698] = 8'h8D;
Memory[19697] = 8'h21;
Memory[19696] = 8'h83;
Memory[19703] = 8'h00;
Memory[19702] = 8'h3B;
Memory[19701] = 8'h2A;
Memory[19700] = 8'h23;
Memory[19707] = 8'h12;
Memory[19706] = 8'h40;
Memory[19705] = 8'h20;
Memory[19704] = 8'h6F;
Memory[19711] = 8'h0B;
Memory[19710] = 8'hCD;
Memory[19709] = 8'h21;
Memory[19708] = 8'h83;
Memory[19715] = 8'h00;
Memory[19714] = 8'h3B;
Memory[19713] = 8'h2A;
Memory[19712] = 8'h23;
Memory[19719] = 8'h12;
Memory[19718] = 8'h40;
Memory[19717] = 8'h20;
Memory[19716] = 8'h6F;
Memory[19723] = 8'h0C;
Memory[19722] = 8'h0D;
Memory[19721] = 8'h21;
Memory[19720] = 8'h83;
Memory[19727] = 8'h00;
Memory[19726] = 8'h3B;
Memory[19725] = 8'h2A;
Memory[19724] = 8'h23;
Memory[19731] = 8'h12;
Memory[19730] = 8'h40;
Memory[19729] = 8'h20;
Memory[19728] = 8'h6F;
Memory[19735] = 8'h0C;
Memory[19734] = 8'h4D;
Memory[19733] = 8'h21;
Memory[19732] = 8'h83;
Memory[19739] = 8'h00;
Memory[19738] = 8'h3B;
Memory[19737] = 8'h2A;
Memory[19736] = 8'h23;
Memory[19743] = 8'h12;
Memory[19742] = 8'h40;
Memory[19741] = 8'h20;
Memory[19740] = 8'h6F;
Memory[19747] = 8'h0C;
Memory[19746] = 8'h8D;
Memory[19745] = 8'h21;
Memory[19744] = 8'h83;
Memory[19751] = 8'h00;
Memory[19750] = 8'h3B;
Memory[19749] = 8'h2A;
Memory[19748] = 8'h23;
Memory[19755] = 8'h12;
Memory[19754] = 8'h40;
Memory[19753] = 8'h20;
Memory[19752] = 8'h6F;
Memory[19759] = 8'h0C;
Memory[19758] = 8'hCD;
Memory[19757] = 8'h21;
Memory[19756] = 8'h83;
Memory[19763] = 8'h00;
Memory[19762] = 8'h3B;
Memory[19761] = 8'h2A;
Memory[19760] = 8'h23;
Memory[19767] = 8'h12;
Memory[19766] = 8'h40;
Memory[19765] = 8'h20;
Memory[19764] = 8'h6F;
Memory[19771] = 8'h0D;
Memory[19770] = 8'h0D;
Memory[19769] = 8'h21;
Memory[19768] = 8'h83;
Memory[19775] = 8'h00;
Memory[19774] = 8'h3B;
Memory[19773] = 8'h2A;
Memory[19772] = 8'h23;
Memory[19779] = 8'h12;
Memory[19778] = 8'h40;
Memory[19777] = 8'h20;
Memory[19776] = 8'h6F;
Memory[19783] = 8'h0D;
Memory[19782] = 8'h4D;
Memory[19781] = 8'h21;
Memory[19780] = 8'h83;
Memory[19787] = 8'h00;
Memory[19786] = 8'h3B;
Memory[19785] = 8'h2A;
Memory[19784] = 8'h23;
Memory[19791] = 8'h12;
Memory[19790] = 8'h40;
Memory[19789] = 8'h20;
Memory[19788] = 8'h6F;
Memory[19795] = 8'h0D;
Memory[19794] = 8'h8D;
Memory[19793] = 8'h21;
Memory[19792] = 8'h83;
Memory[19799] = 8'h00;
Memory[19798] = 8'h3B;
Memory[19797] = 8'h2A;
Memory[19796] = 8'h23;
Memory[19803] = 8'h12;
Memory[19802] = 8'h40;
Memory[19801] = 8'h20;
Memory[19800] = 8'h6F;
Memory[19807] = 8'h0D;
Memory[19806] = 8'hCD;
Memory[19805] = 8'h21;
Memory[19804] = 8'h83;
Memory[19811] = 8'h00;
Memory[19810] = 8'h3B;
Memory[19809] = 8'h2A;
Memory[19808] = 8'h23;
Memory[19815] = 8'h12;
Memory[19814] = 8'h40;
Memory[19813] = 8'h20;
Memory[19812] = 8'h6F;
Memory[19819] = 8'h0E;
Memory[19818] = 8'h0D;
Memory[19817] = 8'h21;
Memory[19816] = 8'h83;
Memory[19823] = 8'h00;
Memory[19822] = 8'h3B;
Memory[19821] = 8'h2A;
Memory[19820] = 8'h23;
Memory[19827] = 8'h12;
Memory[19826] = 8'h40;
Memory[19825] = 8'h20;
Memory[19824] = 8'h6F;
Memory[19831] = 8'h0E;
Memory[19830] = 8'h4D;
Memory[19829] = 8'h21;
Memory[19828] = 8'h83;
Memory[19835] = 8'h00;
Memory[19834] = 8'h3B;
Memory[19833] = 8'h2A;
Memory[19832] = 8'h23;
Memory[19839] = 8'h12;
Memory[19838] = 8'h40;
Memory[19837] = 8'h20;
Memory[19836] = 8'h6F;
Memory[19843] = 8'h0E;
Memory[19842] = 8'h8D;
Memory[19841] = 8'h21;
Memory[19840] = 8'h83;
Memory[19847] = 8'h00;
Memory[19846] = 8'h3B;
Memory[19845] = 8'h2A;
Memory[19844] = 8'h23;
Memory[19851] = 8'h12;
Memory[19850] = 8'h40;
Memory[19849] = 8'h20;
Memory[19848] = 8'h6F;
Memory[19855] = 8'h0E;
Memory[19854] = 8'hCD;
Memory[19853] = 8'h21;
Memory[19852] = 8'h83;
Memory[19859] = 8'h00;
Memory[19858] = 8'h3B;
Memory[19857] = 8'h2A;
Memory[19856] = 8'h23;
Memory[19863] = 8'h12;
Memory[19862] = 8'h40;
Memory[19861] = 8'h20;
Memory[19860] = 8'h6F;
Memory[19867] = 8'h0F;
Memory[19866] = 8'h0D;
Memory[19865] = 8'h21;
Memory[19864] = 8'h83;
Memory[19871] = 8'h00;
Memory[19870] = 8'h3B;
Memory[19869] = 8'h2A;
Memory[19868] = 8'h23;
Memory[19875] = 8'h12;
Memory[19874] = 8'h40;
Memory[19873] = 8'h20;
Memory[19872] = 8'h6F;
Memory[19879] = 8'h0F;
Memory[19878] = 8'h4D;
Memory[19877] = 8'h21;
Memory[19876] = 8'h83;
Memory[19883] = 8'h00;
Memory[19882] = 8'h3B;
Memory[19881] = 8'h2A;
Memory[19880] = 8'h23;
Memory[19887] = 8'h12;
Memory[19886] = 8'h40;
Memory[19885] = 8'h20;
Memory[19884] = 8'h6F;
Memory[19891] = 8'h0F;
Memory[19890] = 8'h8D;
Memory[19889] = 8'h21;
Memory[19888] = 8'h83;
Memory[19895] = 8'h00;
Memory[19894] = 8'h3B;
Memory[19893] = 8'h2A;
Memory[19892] = 8'h23;
Memory[19899] = 8'h12;
Memory[19898] = 8'h40;
Memory[19897] = 8'h20;
Memory[19896] = 8'h6F;
Memory[19903] = 8'h0F;
Memory[19902] = 8'hCD;
Memory[19901] = 8'h21;
Memory[19900] = 8'h83;
Memory[19907] = 8'h00;
Memory[19906] = 8'h3B;
Memory[19905] = 8'h2A;
Memory[19904] = 8'h23;
Memory[19911] = 8'h12;
Memory[19910] = 8'h40;
Memory[19909] = 8'h20;
Memory[19908] = 8'h6F;
Memory[19915] = 8'h10;
Memory[19914] = 8'h0D;
Memory[19913] = 8'h21;
Memory[19912] = 8'h83;
Memory[19919] = 8'h00;
Memory[19918] = 8'h3B;
Memory[19917] = 8'h2A;
Memory[19916] = 8'h23;
Memory[19923] = 8'h12;
Memory[19922] = 8'h40;
Memory[19921] = 8'h20;
Memory[19920] = 8'h6F;
Memory[19927] = 8'h10;
Memory[19926] = 8'h4D;
Memory[19925] = 8'h21;
Memory[19924] = 8'h83;
Memory[19931] = 8'h00;
Memory[19930] = 8'h3B;
Memory[19929] = 8'h2A;
Memory[19928] = 8'h23;
Memory[19935] = 8'h12;
Memory[19934] = 8'h40;
Memory[19933] = 8'h20;
Memory[19932] = 8'h6F;
Memory[19939] = 8'h10;
Memory[19938] = 8'h8D;
Memory[19937] = 8'h21;
Memory[19936] = 8'h83;
Memory[19943] = 8'h00;
Memory[19942] = 8'h3B;
Memory[19941] = 8'h2A;
Memory[19940] = 8'h23;
Memory[19947] = 8'h12;
Memory[19946] = 8'h40;
Memory[19945] = 8'h20;
Memory[19944] = 8'h6F;
Memory[19951] = 8'h10;
Memory[19950] = 8'hCD;
Memory[19949] = 8'h21;
Memory[19948] = 8'h83;
Memory[19955] = 8'h00;
Memory[19954] = 8'h3B;
Memory[19953] = 8'h2A;
Memory[19952] = 8'h23;
Memory[19959] = 8'h12;
Memory[19958] = 8'h40;
Memory[19957] = 8'h20;
Memory[19956] = 8'h6F;
Memory[19963] = 8'h11;
Memory[19962] = 8'h0D;
Memory[19961] = 8'h21;
Memory[19960] = 8'h83;
Memory[19967] = 8'h00;
Memory[19966] = 8'h3B;
Memory[19965] = 8'h2A;
Memory[19964] = 8'h23;
Memory[19971] = 8'h12;
Memory[19970] = 8'h40;
Memory[19969] = 8'h20;
Memory[19968] = 8'h6F;
Memory[19975] = 8'h11;
Memory[19974] = 8'h4D;
Memory[19973] = 8'h21;
Memory[19972] = 8'h83;
Memory[19979] = 8'h00;
Memory[19978] = 8'h3B;
Memory[19977] = 8'h2A;
Memory[19976] = 8'h23;
Memory[19983] = 8'h12;
Memory[19982] = 8'h40;
Memory[19981] = 8'h20;
Memory[19980] = 8'h6F;
Memory[19987] = 8'h11;
Memory[19986] = 8'h8D;
Memory[19985] = 8'h21;
Memory[19984] = 8'h83;
Memory[19991] = 8'h00;
Memory[19990] = 8'h3B;
Memory[19989] = 8'h2A;
Memory[19988] = 8'h23;
Memory[19995] = 8'h12;
Memory[19994] = 8'h40;
Memory[19993] = 8'h20;
Memory[19992] = 8'h6F;
Memory[19999] = 8'h11;
Memory[19998] = 8'hCD;
Memory[19997] = 8'h21;
Memory[19996] = 8'h83;
Memory[20003] = 8'h00;
Memory[20002] = 8'h3B;
Memory[20001] = 8'h2A;
Memory[20000] = 8'h23;
Memory[20007] = 8'h12;
Memory[20006] = 8'h40;
Memory[20005] = 8'h20;
Memory[20004] = 8'h6F;
Memory[20011] = 8'h12;
Memory[20010] = 8'h0D;
Memory[20009] = 8'h21;
Memory[20008] = 8'h83;
Memory[20015] = 8'h00;
Memory[20014] = 8'h3B;
Memory[20013] = 8'h2A;
Memory[20012] = 8'h23;
Memory[20019] = 8'h12;
Memory[20018] = 8'h40;
Memory[20017] = 8'h20;
Memory[20016] = 8'h6F;
Memory[20023] = 8'h12;
Memory[20022] = 8'h4D;
Memory[20021] = 8'h21;
Memory[20020] = 8'h83;
Memory[20027] = 8'h00;
Memory[20026] = 8'h3B;
Memory[20025] = 8'h2A;
Memory[20024] = 8'h23;
Memory[20031] = 8'h12;
Memory[20030] = 8'h40;
Memory[20029] = 8'h20;
Memory[20028] = 8'h6F;
Memory[20035] = 8'h12;
Memory[20034] = 8'h8D;
Memory[20033] = 8'h21;
Memory[20032] = 8'h83;
Memory[20039] = 8'h00;
Memory[20038] = 8'h3B;
Memory[20037] = 8'h2A;
Memory[20036] = 8'h23;
Memory[20043] = 8'h12;
Memory[20042] = 8'h40;
Memory[20041] = 8'h20;
Memory[20040] = 8'h6F;
Memory[20047] = 8'h12;
Memory[20046] = 8'hCD;
Memory[20045] = 8'h21;
Memory[20044] = 8'h83;
Memory[20051] = 8'h00;
Memory[20050] = 8'h3B;
Memory[20049] = 8'h2A;
Memory[20048] = 8'h23;
Memory[20055] = 8'h12;
Memory[20054] = 8'h40;
Memory[20053] = 8'h20;
Memory[20052] = 8'h6F;
Memory[20059] = 8'h13;
Memory[20058] = 8'h0D;
Memory[20057] = 8'h21;
Memory[20056] = 8'h83;
Memory[20063] = 8'h00;
Memory[20062] = 8'h3B;
Memory[20061] = 8'h2A;
Memory[20060] = 8'h23;
Memory[20067] = 8'h12;
Memory[20066] = 8'h40;
Memory[20065] = 8'h20;
Memory[20064] = 8'h6F;
Memory[20071] = 8'h13;
Memory[20070] = 8'h4D;
Memory[20069] = 8'h21;
Memory[20068] = 8'h83;
Memory[20075] = 8'h00;
Memory[20074] = 8'h3B;
Memory[20073] = 8'h2A;
Memory[20072] = 8'h23;
Memory[20079] = 8'h12;
Memory[20078] = 8'h40;
Memory[20077] = 8'h20;
Memory[20076] = 8'h6F;
Memory[20083] = 8'h13;
Memory[20082] = 8'h8D;
Memory[20081] = 8'h21;
Memory[20080] = 8'h83;
Memory[20087] = 8'h00;
Memory[20086] = 8'h3B;
Memory[20085] = 8'h2A;
Memory[20084] = 8'h23;
Memory[20091] = 8'h12;
Memory[20090] = 8'h40;
Memory[20089] = 8'h20;
Memory[20088] = 8'h6F;
Memory[20095] = 8'h13;
Memory[20094] = 8'hCD;
Memory[20093] = 8'h21;
Memory[20092] = 8'h83;
Memory[20099] = 8'h00;
Memory[20098] = 8'h3B;
Memory[20097] = 8'h2A;
Memory[20096] = 8'h23;
Memory[20103] = 8'h12;
Memory[20102] = 8'h40;
Memory[20101] = 8'h20;
Memory[20100] = 8'h6F;
Memory[20107] = 8'h14;
Memory[20106] = 8'h0D;
Memory[20105] = 8'h21;
Memory[20104] = 8'h83;
Memory[20111] = 8'h00;
Memory[20110] = 8'h3B;
Memory[20109] = 8'h2A;
Memory[20108] = 8'h23;
Memory[20115] = 8'h12;
Memory[20114] = 8'h40;
Memory[20113] = 8'h20;
Memory[20112] = 8'h6F;
Memory[20119] = 8'h14;
Memory[20118] = 8'h4D;
Memory[20117] = 8'h21;
Memory[20116] = 8'h83;
Memory[20123] = 8'h00;
Memory[20122] = 8'h3B;
Memory[20121] = 8'h2A;
Memory[20120] = 8'h23;
Memory[20127] = 8'h12;
Memory[20126] = 8'h40;
Memory[20125] = 8'h20;
Memory[20124] = 8'h6F;
Memory[20131] = 8'h14;
Memory[20130] = 8'h8D;
Memory[20129] = 8'h21;
Memory[20128] = 8'h83;
Memory[20135] = 8'h00;
Memory[20134] = 8'h3B;
Memory[20133] = 8'h2A;
Memory[20132] = 8'h23;
Memory[20139] = 8'h12;
Memory[20138] = 8'h40;
Memory[20137] = 8'h20;
Memory[20136] = 8'h6F;
Memory[20143] = 8'h14;
Memory[20142] = 8'hCD;
Memory[20141] = 8'h21;
Memory[20140] = 8'h83;
Memory[20147] = 8'h00;
Memory[20146] = 8'h3B;
Memory[20145] = 8'h2A;
Memory[20144] = 8'h23;
Memory[20151] = 8'h12;
Memory[20150] = 8'h40;
Memory[20149] = 8'h20;
Memory[20148] = 8'h6F;
Memory[20155] = 8'h15;
Memory[20154] = 8'h0D;
Memory[20153] = 8'h21;
Memory[20152] = 8'h83;
Memory[20159] = 8'h00;
Memory[20158] = 8'h3B;
Memory[20157] = 8'h2A;
Memory[20156] = 8'h23;
Memory[20163] = 8'h12;
Memory[20162] = 8'h40;
Memory[20161] = 8'h20;
Memory[20160] = 8'h6F;
Memory[20167] = 8'h15;
Memory[20166] = 8'h4D;
Memory[20165] = 8'h21;
Memory[20164] = 8'h83;
Memory[20171] = 8'h00;
Memory[20170] = 8'h3B;
Memory[20169] = 8'h2A;
Memory[20168] = 8'h23;
Memory[20175] = 8'h12;
Memory[20174] = 8'h40;
Memory[20173] = 8'h20;
Memory[20172] = 8'h6F;
Memory[20179] = 8'h15;
Memory[20178] = 8'h8D;
Memory[20177] = 8'h21;
Memory[20176] = 8'h83;
Memory[20183] = 8'h00;
Memory[20182] = 8'h3B;
Memory[20181] = 8'h2A;
Memory[20180] = 8'h23;
Memory[20187] = 8'h12;
Memory[20186] = 8'h40;
Memory[20185] = 8'h20;
Memory[20184] = 8'h6F;
Memory[20191] = 8'h15;
Memory[20190] = 8'hCD;
Memory[20189] = 8'h21;
Memory[20188] = 8'h83;
Memory[20195] = 8'h00;
Memory[20194] = 8'h3B;
Memory[20193] = 8'h2A;
Memory[20192] = 8'h23;
Memory[20199] = 8'h12;
Memory[20198] = 8'h40;
Memory[20197] = 8'h20;
Memory[20196] = 8'h6F;
Memory[20203] = 8'h16;
Memory[20202] = 8'h0D;
Memory[20201] = 8'h21;
Memory[20200] = 8'h83;
Memory[20207] = 8'h00;
Memory[20206] = 8'h3B;
Memory[20205] = 8'h2A;
Memory[20204] = 8'h23;
Memory[20211] = 8'h12;
Memory[20210] = 8'h40;
Memory[20209] = 8'h20;
Memory[20208] = 8'h6F;
Memory[20215] = 8'h16;
Memory[20214] = 8'h4D;
Memory[20213] = 8'h21;
Memory[20212] = 8'h83;
Memory[20219] = 8'h00;
Memory[20218] = 8'h3B;
Memory[20217] = 8'h2A;
Memory[20216] = 8'h23;
Memory[20223] = 8'h12;
Memory[20222] = 8'h40;
Memory[20221] = 8'h20;
Memory[20220] = 8'h6F;
Memory[20227] = 8'h16;
Memory[20226] = 8'h8D;
Memory[20225] = 8'h21;
Memory[20224] = 8'h83;
Memory[20231] = 8'h00;
Memory[20230] = 8'h3B;
Memory[20229] = 8'h2A;
Memory[20228] = 8'h23;
Memory[20235] = 8'h12;
Memory[20234] = 8'h40;
Memory[20233] = 8'h20;
Memory[20232] = 8'h6F;
Memory[20239] = 8'h16;
Memory[20238] = 8'hCD;
Memory[20237] = 8'h21;
Memory[20236] = 8'h83;
Memory[20243] = 8'h00;
Memory[20242] = 8'h3B;
Memory[20241] = 8'h2A;
Memory[20240] = 8'h23;
Memory[20247] = 8'h12;
Memory[20246] = 8'h40;
Memory[20245] = 8'h20;
Memory[20244] = 8'h6F;
Memory[20251] = 8'h17;
Memory[20250] = 8'h0D;
Memory[20249] = 8'h21;
Memory[20248] = 8'h83;
Memory[20255] = 8'h00;
Memory[20254] = 8'h3B;
Memory[20253] = 8'h2A;
Memory[20252] = 8'h23;
Memory[20259] = 8'h12;
Memory[20258] = 8'h40;
Memory[20257] = 8'h20;
Memory[20256] = 8'h6F;
Memory[20263] = 8'h17;
Memory[20262] = 8'h4D;
Memory[20261] = 8'h21;
Memory[20260] = 8'h83;
Memory[20267] = 8'h00;
Memory[20266] = 8'h3B;
Memory[20265] = 8'h2A;
Memory[20264] = 8'h23;
Memory[20271] = 8'h12;
Memory[20270] = 8'h40;
Memory[20269] = 8'h20;
Memory[20268] = 8'h6F;
Memory[20275] = 8'h17;
Memory[20274] = 8'h8D;
Memory[20273] = 8'h21;
Memory[20272] = 8'h83;
Memory[20279] = 8'h00;
Memory[20278] = 8'h3B;
Memory[20277] = 8'h2A;
Memory[20276] = 8'h23;
Memory[20283] = 8'h12;
Memory[20282] = 8'h40;
Memory[20281] = 8'h20;
Memory[20280] = 8'h6F;
Memory[20287] = 8'h17;
Memory[20286] = 8'hCD;
Memory[20285] = 8'h21;
Memory[20284] = 8'h83;
Memory[20291] = 8'h00;
Memory[20290] = 8'h3B;
Memory[20289] = 8'h2A;
Memory[20288] = 8'h23;
Memory[20295] = 8'h12;
Memory[20294] = 8'h40;
Memory[20293] = 8'h20;
Memory[20292] = 8'h6F;
Memory[20299] = 8'h18;
Memory[20298] = 8'h0D;
Memory[20297] = 8'h21;
Memory[20296] = 8'h83;
Memory[20303] = 8'h00;
Memory[20302] = 8'h3B;
Memory[20301] = 8'h2A;
Memory[20300] = 8'h23;
Memory[20307] = 8'h12;
Memory[20306] = 8'h40;
Memory[20305] = 8'h20;
Memory[20304] = 8'h6F;
Memory[20311] = 8'h18;
Memory[20310] = 8'h4D;
Memory[20309] = 8'h21;
Memory[20308] = 8'h83;
Memory[20315] = 8'h00;
Memory[20314] = 8'h3B;
Memory[20313] = 8'h2A;
Memory[20312] = 8'h23;
Memory[20319] = 8'h12;
Memory[20318] = 8'h40;
Memory[20317] = 8'h20;
Memory[20316] = 8'h6F;
Memory[20323] = 8'h18;
Memory[20322] = 8'h8D;
Memory[20321] = 8'h21;
Memory[20320] = 8'h83;
Memory[20327] = 8'h00;
Memory[20326] = 8'h3B;
Memory[20325] = 8'h2A;
Memory[20324] = 8'h23;
Memory[20331] = 8'h12;
Memory[20330] = 8'h40;
Memory[20329] = 8'h20;
Memory[20328] = 8'h6F;
Memory[20335] = 8'h18;
Memory[20334] = 8'hCD;
Memory[20333] = 8'h21;
Memory[20332] = 8'h83;
Memory[20339] = 8'h00;
Memory[20338] = 8'h3B;
Memory[20337] = 8'h2A;
Memory[20336] = 8'h23;
Memory[20343] = 8'h12;
Memory[20342] = 8'h40;
Memory[20341] = 8'h20;
Memory[20340] = 8'h6F;
Memory[20347] = 8'h19;
Memory[20346] = 8'h0D;
Memory[20345] = 8'h21;
Memory[20344] = 8'h83;
Memory[20351] = 8'h00;
Memory[20350] = 8'h3B;
Memory[20349] = 8'h2A;
Memory[20348] = 8'h23;
Memory[20355] = 8'h12;
Memory[20354] = 8'h40;
Memory[20353] = 8'h20;
Memory[20352] = 8'h6F;
Memory[20359] = 8'h19;
Memory[20358] = 8'h4D;
Memory[20357] = 8'h21;
Memory[20356] = 8'h83;
Memory[20363] = 8'h00;
Memory[20362] = 8'h3B;
Memory[20361] = 8'h2A;
Memory[20360] = 8'h23;
Memory[20367] = 8'h12;
Memory[20366] = 8'h40;
Memory[20365] = 8'h20;
Memory[20364] = 8'h6F;
Memory[20371] = 8'h19;
Memory[20370] = 8'h8D;
Memory[20369] = 8'h21;
Memory[20368] = 8'h83;
Memory[20375] = 8'h00;
Memory[20374] = 8'h3B;
Memory[20373] = 8'h2A;
Memory[20372] = 8'h23;
Memory[20379] = 8'h12;
Memory[20378] = 8'h40;
Memory[20377] = 8'h20;
Memory[20376] = 8'h6F;
Memory[20383] = 8'h19;
Memory[20382] = 8'hCD;
Memory[20381] = 8'h21;
Memory[20380] = 8'h83;
Memory[20387] = 8'h00;
Memory[20386] = 8'h3B;
Memory[20385] = 8'h2A;
Memory[20384] = 8'h23;
Memory[20391] = 8'h12;
Memory[20390] = 8'h40;
Memory[20389] = 8'h20;
Memory[20388] = 8'h6F;
Memory[20395] = 8'h1A;
Memory[20394] = 8'h0D;
Memory[20393] = 8'h21;
Memory[20392] = 8'h83;
Memory[20399] = 8'h00;
Memory[20398] = 8'h3B;
Memory[20397] = 8'h2A;
Memory[20396] = 8'h23;
Memory[20403] = 8'h12;
Memory[20402] = 8'h40;
Memory[20401] = 8'h20;
Memory[20400] = 8'h6F;
Memory[20407] = 8'h1A;
Memory[20406] = 8'h4D;
Memory[20405] = 8'h21;
Memory[20404] = 8'h83;
Memory[20411] = 8'h00;
Memory[20410] = 8'h3B;
Memory[20409] = 8'h2A;
Memory[20408] = 8'h23;
Memory[20415] = 8'h12;
Memory[20414] = 8'h40;
Memory[20413] = 8'h20;
Memory[20412] = 8'h6F;
Memory[20419] = 8'h1A;
Memory[20418] = 8'h8D;
Memory[20417] = 8'h21;
Memory[20416] = 8'h83;
Memory[20423] = 8'h00;
Memory[20422] = 8'h3B;
Memory[20421] = 8'h2A;
Memory[20420] = 8'h23;
Memory[20427] = 8'h12;
Memory[20426] = 8'h40;
Memory[20425] = 8'h20;
Memory[20424] = 8'h6F;
Memory[20431] = 8'h1A;
Memory[20430] = 8'hCD;
Memory[20429] = 8'h21;
Memory[20428] = 8'h83;
Memory[20435] = 8'h00;
Memory[20434] = 8'h3B;
Memory[20433] = 8'h2A;
Memory[20432] = 8'h23;
Memory[20439] = 8'h12;
Memory[20438] = 8'h40;
Memory[20437] = 8'h20;
Memory[20436] = 8'h6F;
Memory[20443] = 8'h1B;
Memory[20442] = 8'h0D;
Memory[20441] = 8'h21;
Memory[20440] = 8'h83;
Memory[20447] = 8'h00;
Memory[20446] = 8'h3B;
Memory[20445] = 8'h2A;
Memory[20444] = 8'h23;
Memory[20451] = 8'h12;
Memory[20450] = 8'h40;
Memory[20449] = 8'h20;
Memory[20448] = 8'h6F;
Memory[20455] = 8'h1B;
Memory[20454] = 8'h4D;
Memory[20453] = 8'h21;
Memory[20452] = 8'h83;
Memory[20459] = 8'h00;
Memory[20458] = 8'h3B;
Memory[20457] = 8'h2A;
Memory[20456] = 8'h23;
Memory[20463] = 8'h12;
Memory[20462] = 8'h40;
Memory[20461] = 8'h20;
Memory[20460] = 8'h6F;
Memory[20467] = 8'h1B;
Memory[20466] = 8'h8D;
Memory[20465] = 8'h21;
Memory[20464] = 8'h83;
Memory[20471] = 8'h00;
Memory[20470] = 8'h3B;
Memory[20469] = 8'h2A;
Memory[20468] = 8'h23;
Memory[20475] = 8'h12;
Memory[20474] = 8'h40;
Memory[20473] = 8'h20;
Memory[20472] = 8'h6F;
Memory[20479] = 8'h1B;
Memory[20478] = 8'hCD;
Memory[20477] = 8'h21;
Memory[20476] = 8'h83;
Memory[20483] = 8'h00;
Memory[20482] = 8'h3B;
Memory[20481] = 8'h2A;
Memory[20480] = 8'h23;
Memory[20487] = 8'h12;
Memory[20486] = 8'h40;
Memory[20485] = 8'h20;
Memory[20484] = 8'h6F;
Memory[20491] = 8'h1C;
Memory[20490] = 8'h0D;
Memory[20489] = 8'h21;
Memory[20488] = 8'h83;
Memory[20495] = 8'h00;
Memory[20494] = 8'h3B;
Memory[20493] = 8'h2A;
Memory[20492] = 8'h23;
Memory[20499] = 8'h12;
Memory[20498] = 8'h40;
Memory[20497] = 8'h20;
Memory[20496] = 8'h6F;
Memory[20503] = 8'h1C;
Memory[20502] = 8'h4D;
Memory[20501] = 8'h21;
Memory[20500] = 8'h83;
Memory[20507] = 8'h00;
Memory[20506] = 8'h3B;
Memory[20505] = 8'h2A;
Memory[20504] = 8'h23;
Memory[20511] = 8'h12;
Memory[20510] = 8'h40;
Memory[20509] = 8'h20;
Memory[20508] = 8'h6F;
Memory[20515] = 8'h1C;
Memory[20514] = 8'h8D;
Memory[20513] = 8'h21;
Memory[20512] = 8'h83;
Memory[20519] = 8'h00;
Memory[20518] = 8'h3B;
Memory[20517] = 8'h2A;
Memory[20516] = 8'h23;
Memory[20523] = 8'h12;
Memory[20522] = 8'h40;
Memory[20521] = 8'h20;
Memory[20520] = 8'h6F;
Memory[20527] = 8'h1C;
Memory[20526] = 8'hCD;
Memory[20525] = 8'h21;
Memory[20524] = 8'h83;
Memory[20531] = 8'h00;
Memory[20530] = 8'h3B;
Memory[20529] = 8'h2A;
Memory[20528] = 8'h23;
Memory[20535] = 8'h12;
Memory[20534] = 8'h40;
Memory[20533] = 8'h20;
Memory[20532] = 8'h6F;
Memory[20539] = 8'h1D;
Memory[20538] = 8'h0D;
Memory[20537] = 8'h21;
Memory[20536] = 8'h83;
Memory[20543] = 8'h00;
Memory[20542] = 8'h3B;
Memory[20541] = 8'h2A;
Memory[20540] = 8'h23;
Memory[20547] = 8'h12;
Memory[20546] = 8'h40;
Memory[20545] = 8'h20;
Memory[20544] = 8'h6F;
Memory[20551] = 8'h1D;
Memory[20550] = 8'h4D;
Memory[20549] = 8'h21;
Memory[20548] = 8'h83;
Memory[20555] = 8'h00;
Memory[20554] = 8'h3B;
Memory[20553] = 8'h2A;
Memory[20552] = 8'h23;
Memory[20559] = 8'h12;
Memory[20558] = 8'h40;
Memory[20557] = 8'h20;
Memory[20556] = 8'h6F;
Memory[20563] = 8'h1D;
Memory[20562] = 8'h8D;
Memory[20561] = 8'h21;
Memory[20560] = 8'h83;
Memory[20567] = 8'h00;
Memory[20566] = 8'h3B;
Memory[20565] = 8'h2A;
Memory[20564] = 8'h23;
Memory[20571] = 8'h12;
Memory[20570] = 8'h40;
Memory[20569] = 8'h20;
Memory[20568] = 8'h6F;
Memory[20575] = 8'h1D;
Memory[20574] = 8'hCD;
Memory[20573] = 8'h21;
Memory[20572] = 8'h83;
Memory[20579] = 8'h00;
Memory[20578] = 8'h3B;
Memory[20577] = 8'h2A;
Memory[20576] = 8'h23;
Memory[20583] = 8'h12;
Memory[20582] = 8'h40;
Memory[20581] = 8'h20;
Memory[20580] = 8'h6F;
Memory[20587] = 8'h1E;
Memory[20586] = 8'h0D;
Memory[20585] = 8'h21;
Memory[20584] = 8'h83;
Memory[20591] = 8'h00;
Memory[20590] = 8'h3B;
Memory[20589] = 8'h2A;
Memory[20588] = 8'h23;
Memory[20595] = 8'h12;
Memory[20594] = 8'h40;
Memory[20593] = 8'h20;
Memory[20592] = 8'h6F;
Memory[20599] = 8'h1E;
Memory[20598] = 8'h4D;
Memory[20597] = 8'h21;
Memory[20596] = 8'h83;
Memory[20603] = 8'h00;
Memory[20602] = 8'h3B;
Memory[20601] = 8'h2A;
Memory[20600] = 8'h23;
Memory[20607] = 8'h12;
Memory[20606] = 8'h40;
Memory[20605] = 8'h20;
Memory[20604] = 8'h6F;
Memory[20611] = 8'h1E;
Memory[20610] = 8'h8D;
Memory[20609] = 8'h21;
Memory[20608] = 8'h83;
Memory[20615] = 8'h00;
Memory[20614] = 8'h3B;
Memory[20613] = 8'h2A;
Memory[20612] = 8'h23;
Memory[20619] = 8'h12;
Memory[20618] = 8'h40;
Memory[20617] = 8'h20;
Memory[20616] = 8'h6F;
Memory[20623] = 8'h1E;
Memory[20622] = 8'hCD;
Memory[20621] = 8'h21;
Memory[20620] = 8'h83;
Memory[20627] = 8'h00;
Memory[20626] = 8'h3B;
Memory[20625] = 8'h2A;
Memory[20624] = 8'h23;
Memory[20631] = 8'h12;
Memory[20630] = 8'h40;
Memory[20629] = 8'h20;
Memory[20628] = 8'h6F;
Memory[20635] = 8'h1F;
Memory[20634] = 8'h0D;
Memory[20633] = 8'h21;
Memory[20632] = 8'h83;
Memory[20639] = 8'h00;
Memory[20638] = 8'h3B;
Memory[20637] = 8'h2A;
Memory[20636] = 8'h23;
Memory[20643] = 8'h12;
Memory[20642] = 8'h40;
Memory[20641] = 8'h20;
Memory[20640] = 8'h6F;
Memory[20647] = 8'h1F;
Memory[20646] = 8'h4D;
Memory[20645] = 8'h21;
Memory[20644] = 8'h83;
Memory[20651] = 8'h00;
Memory[20650] = 8'h3B;
Memory[20649] = 8'h2A;
Memory[20648] = 8'h23;
Memory[20655] = 8'h12;
Memory[20654] = 8'h40;
Memory[20653] = 8'h20;
Memory[20652] = 8'h6F;
Memory[20659] = 8'h1F;
Memory[20658] = 8'h8D;
Memory[20657] = 8'h21;
Memory[20656] = 8'h83;
Memory[20663] = 8'h00;
Memory[20662] = 8'h3B;
Memory[20661] = 8'h2A;
Memory[20660] = 8'h23;
Memory[20667] = 8'h12;
Memory[20666] = 8'h40;
Memory[20665] = 8'h20;
Memory[20664] = 8'h6F;
Memory[20671] = 8'h1F;
Memory[20670] = 8'hCD;
Memory[20669] = 8'h21;
Memory[20668] = 8'h83;
Memory[20675] = 8'h00;
Memory[20674] = 8'h3B;
Memory[20673] = 8'h2A;
Memory[20672] = 8'h23;
Memory[20679] = 8'h12;
Memory[20678] = 8'h40;
Memory[20677] = 8'h20;
Memory[20676] = 8'h6F;
Memory[20683] = 8'h20;
Memory[20682] = 8'h0D;
Memory[20681] = 8'h21;
Memory[20680] = 8'h83;
Memory[20687] = 8'h00;
Memory[20686] = 8'h3B;
Memory[20685] = 8'h2A;
Memory[20684] = 8'h23;
Memory[20691] = 8'h12;
Memory[20690] = 8'h40;
Memory[20689] = 8'h20;
Memory[20688] = 8'h6F;
Memory[20695] = 8'h20;
Memory[20694] = 8'h4D;
Memory[20693] = 8'h21;
Memory[20692] = 8'h83;
Memory[20699] = 8'h00;
Memory[20698] = 8'h3B;
Memory[20697] = 8'h2A;
Memory[20696] = 8'h23;
Memory[20703] = 8'h12;
Memory[20702] = 8'h40;
Memory[20701] = 8'h20;
Memory[20700] = 8'h6F;
Memory[20707] = 8'h20;
Memory[20706] = 8'h8D;
Memory[20705] = 8'h21;
Memory[20704] = 8'h83;
Memory[20711] = 8'h00;
Memory[20710] = 8'h3B;
Memory[20709] = 8'h2A;
Memory[20708] = 8'h23;
Memory[20715] = 8'h12;
Memory[20714] = 8'h40;
Memory[20713] = 8'h20;
Memory[20712] = 8'h6F;
Memory[20719] = 8'h20;
Memory[20718] = 8'hCD;
Memory[20717] = 8'h21;
Memory[20716] = 8'h83;
Memory[20723] = 8'h00;
Memory[20722] = 8'h3B;
Memory[20721] = 8'h2A;
Memory[20720] = 8'h23;
Memory[20727] = 8'h12;
Memory[20726] = 8'h40;
Memory[20725] = 8'h20;
Memory[20724] = 8'h6F;
Memory[20731] = 8'h21;
Memory[20730] = 8'h0D;
Memory[20729] = 8'h21;
Memory[20728] = 8'h83;
Memory[20735] = 8'h00;
Memory[20734] = 8'h3B;
Memory[20733] = 8'h2A;
Memory[20732] = 8'h23;
Memory[20739] = 8'h12;
Memory[20738] = 8'h40;
Memory[20737] = 8'h20;
Memory[20736] = 8'h6F;
Memory[20743] = 8'h21;
Memory[20742] = 8'h4D;
Memory[20741] = 8'h21;
Memory[20740] = 8'h83;
Memory[20747] = 8'h00;
Memory[20746] = 8'h3B;
Memory[20745] = 8'h2A;
Memory[20744] = 8'h23;
Memory[20751] = 8'h12;
Memory[20750] = 8'h40;
Memory[20749] = 8'h20;
Memory[20748] = 8'h6F;
Memory[20755] = 8'h21;
Memory[20754] = 8'h8D;
Memory[20753] = 8'h21;
Memory[20752] = 8'h83;
Memory[20759] = 8'h00;
Memory[20758] = 8'h3B;
Memory[20757] = 8'h2A;
Memory[20756] = 8'h23;
Memory[20763] = 8'h12;
Memory[20762] = 8'h40;
Memory[20761] = 8'h20;
Memory[20760] = 8'h6F;
Memory[20767] = 8'h21;
Memory[20766] = 8'hCD;
Memory[20765] = 8'h21;
Memory[20764] = 8'h83;
Memory[20771] = 8'h00;
Memory[20770] = 8'h3B;
Memory[20769] = 8'h2A;
Memory[20768] = 8'h23;
Memory[20775] = 8'h12;
Memory[20774] = 8'h40;
Memory[20773] = 8'h20;
Memory[20772] = 8'h6F;
Memory[20779] = 8'h22;
Memory[20778] = 8'h0D;
Memory[20777] = 8'h21;
Memory[20776] = 8'h83;
Memory[20783] = 8'h00;
Memory[20782] = 8'h3B;
Memory[20781] = 8'h2A;
Memory[20780] = 8'h23;
Memory[20787] = 8'h12;
Memory[20786] = 8'h40;
Memory[20785] = 8'h20;
Memory[20784] = 8'h6F;
Memory[20791] = 8'h22;
Memory[20790] = 8'h4D;
Memory[20789] = 8'h21;
Memory[20788] = 8'h83;
Memory[20795] = 8'h00;
Memory[20794] = 8'h3B;
Memory[20793] = 8'h2A;
Memory[20792] = 8'h23;
Memory[20799] = 8'h12;
Memory[20798] = 8'h40;
Memory[20797] = 8'h20;
Memory[20796] = 8'h6F;
Memory[20803] = 8'h22;
Memory[20802] = 8'h8D;
Memory[20801] = 8'h21;
Memory[20800] = 8'h83;
Memory[20807] = 8'h00;
Memory[20806] = 8'h3B;
Memory[20805] = 8'h2A;
Memory[20804] = 8'h23;
Memory[20811] = 8'h12;
Memory[20810] = 8'h40;
Memory[20809] = 8'h20;
Memory[20808] = 8'h6F;
Memory[20815] = 8'h22;
Memory[20814] = 8'hCD;
Memory[20813] = 8'h21;
Memory[20812] = 8'h83;
Memory[20819] = 8'h00;
Memory[20818] = 8'h3B;
Memory[20817] = 8'h2A;
Memory[20816] = 8'h23;
Memory[20823] = 8'h12;
Memory[20822] = 8'h40;
Memory[20821] = 8'h20;
Memory[20820] = 8'h6F;
Memory[20827] = 8'h23;
Memory[20826] = 8'h0D;
Memory[20825] = 8'h21;
Memory[20824] = 8'h83;
Memory[20831] = 8'h00;
Memory[20830] = 8'h3B;
Memory[20829] = 8'h2A;
Memory[20828] = 8'h23;
Memory[20835] = 8'h12;
Memory[20834] = 8'h40;
Memory[20833] = 8'h20;
Memory[20832] = 8'h6F;
Memory[20839] = 8'h23;
Memory[20838] = 8'h4D;
Memory[20837] = 8'h21;
Memory[20836] = 8'h83;
Memory[20843] = 8'h00;
Memory[20842] = 8'h3B;
Memory[20841] = 8'h2A;
Memory[20840] = 8'h23;
Memory[20847] = 8'h12;
Memory[20846] = 8'h40;
Memory[20845] = 8'h20;
Memory[20844] = 8'h6F;
Memory[20851] = 8'h23;
Memory[20850] = 8'h8D;
Memory[20849] = 8'h21;
Memory[20848] = 8'h83;
Memory[20855] = 8'h00;
Memory[20854] = 8'h3B;
Memory[20853] = 8'h2A;
Memory[20852] = 8'h23;
Memory[20859] = 8'h12;
Memory[20858] = 8'h40;
Memory[20857] = 8'h20;
Memory[20856] = 8'h6F;
Memory[20863] = 8'h23;
Memory[20862] = 8'hCD;
Memory[20861] = 8'h21;
Memory[20860] = 8'h83;
Memory[20867] = 8'h00;
Memory[20866] = 8'h3B;
Memory[20865] = 8'h2A;
Memory[20864] = 8'h23;
Memory[20871] = 8'h12;
Memory[20870] = 8'h40;
Memory[20869] = 8'h20;
Memory[20868] = 8'h6F;
Memory[20875] = 8'h24;
Memory[20874] = 8'h0D;
Memory[20873] = 8'h21;
Memory[20872] = 8'h83;
Memory[20879] = 8'h00;
Memory[20878] = 8'h3B;
Memory[20877] = 8'h2A;
Memory[20876] = 8'h23;
Memory[20883] = 8'h12;
Memory[20882] = 8'h40;
Memory[20881] = 8'h20;
Memory[20880] = 8'h6F;
Memory[20887] = 8'h24;
Memory[20886] = 8'h4D;
Memory[20885] = 8'h21;
Memory[20884] = 8'h83;
Memory[20891] = 8'h00;
Memory[20890] = 8'h3B;
Memory[20889] = 8'h2A;
Memory[20888] = 8'h23;
Memory[20895] = 8'h12;
Memory[20894] = 8'h40;
Memory[20893] = 8'h20;
Memory[20892] = 8'h6F;
Memory[20899] = 8'h24;
Memory[20898] = 8'h8D;
Memory[20897] = 8'h21;
Memory[20896] = 8'h83;
Memory[20903] = 8'h00;
Memory[20902] = 8'h3B;
Memory[20901] = 8'h2A;
Memory[20900] = 8'h23;
Memory[20907] = 8'h12;
Memory[20906] = 8'h40;
Memory[20905] = 8'h20;
Memory[20904] = 8'h6F;
Memory[20911] = 8'h24;
Memory[20910] = 8'hCD;
Memory[20909] = 8'h21;
Memory[20908] = 8'h83;
Memory[20915] = 8'h00;
Memory[20914] = 8'h3B;
Memory[20913] = 8'h2A;
Memory[20912] = 8'h23;
Memory[20919] = 8'h12;
Memory[20918] = 8'h40;
Memory[20917] = 8'h20;
Memory[20916] = 8'h6F;
Memory[20923] = 8'h25;
Memory[20922] = 8'h0D;
Memory[20921] = 8'h21;
Memory[20920] = 8'h83;
Memory[20927] = 8'h00;
Memory[20926] = 8'h3B;
Memory[20925] = 8'h2A;
Memory[20924] = 8'h23;
Memory[20931] = 8'h12;
Memory[20930] = 8'h40;
Memory[20929] = 8'h20;
Memory[20928] = 8'h6F;
Memory[20935] = 8'h25;
Memory[20934] = 8'h4D;
Memory[20933] = 8'h21;
Memory[20932] = 8'h83;
Memory[20939] = 8'h00;
Memory[20938] = 8'h3B;
Memory[20937] = 8'h2A;
Memory[20936] = 8'h23;
Memory[20943] = 8'h12;
Memory[20942] = 8'h40;
Memory[20941] = 8'h20;
Memory[20940] = 8'h6F;
Memory[20947] = 8'h25;
Memory[20946] = 8'h8D;
Memory[20945] = 8'h21;
Memory[20944] = 8'h83;
Memory[20951] = 8'h00;
Memory[20950] = 8'h3B;
Memory[20949] = 8'h2A;
Memory[20948] = 8'h23;
Memory[20955] = 8'h12;
Memory[20954] = 8'h40;
Memory[20953] = 8'h20;
Memory[20952] = 8'h6F;
Memory[20959] = 8'h25;
Memory[20958] = 8'hCD;
Memory[20957] = 8'h21;
Memory[20956] = 8'h83;
Memory[20963] = 8'h00;
Memory[20962] = 8'h3B;
Memory[20961] = 8'h2A;
Memory[20960] = 8'h23;
Memory[20967] = 8'h12;
Memory[20966] = 8'h40;
Memory[20965] = 8'h20;
Memory[20964] = 8'h6F;
Memory[20971] = 8'h26;
Memory[20970] = 8'h0D;
Memory[20969] = 8'h21;
Memory[20968] = 8'h83;
Memory[20975] = 8'h00;
Memory[20974] = 8'h3B;
Memory[20973] = 8'h2A;
Memory[20972] = 8'h23;
Memory[20979] = 8'h12;
Memory[20978] = 8'h40;
Memory[20977] = 8'h20;
Memory[20976] = 8'h6F;
Memory[20983] = 8'h26;
Memory[20982] = 8'h4D;
Memory[20981] = 8'h21;
Memory[20980] = 8'h83;
Memory[20987] = 8'h00;
Memory[20986] = 8'h3B;
Memory[20985] = 8'h2A;
Memory[20984] = 8'h23;
Memory[20991] = 8'h12;
Memory[20990] = 8'h40;
Memory[20989] = 8'h20;
Memory[20988] = 8'h6F;
Memory[20995] = 8'h26;
Memory[20994] = 8'h8D;
Memory[20993] = 8'h21;
Memory[20992] = 8'h83;
Memory[20999] = 8'h00;
Memory[20998] = 8'h3B;
Memory[20997] = 8'h2A;
Memory[20996] = 8'h23;
Memory[21003] = 8'h12;
Memory[21002] = 8'h40;
Memory[21001] = 8'h20;
Memory[21000] = 8'h6F;
Memory[21007] = 8'h26;
Memory[21006] = 8'hCD;
Memory[21005] = 8'h21;
Memory[21004] = 8'h83;
Memory[21011] = 8'h00;
Memory[21010] = 8'h3B;
Memory[21009] = 8'h2A;
Memory[21008] = 8'h23;
Memory[21015] = 8'h12;
Memory[21014] = 8'h40;
Memory[21013] = 8'h20;
Memory[21012] = 8'h6F;
Memory[21019] = 8'h27;
Memory[21018] = 8'h0D;
Memory[21017] = 8'h21;
Memory[21016] = 8'h83;
Memory[21023] = 8'h00;
Memory[21022] = 8'h3B;
Memory[21021] = 8'h2A;
Memory[21020] = 8'h23;
Memory[21027] = 8'h12;
Memory[21026] = 8'h40;
Memory[21025] = 8'h20;
Memory[21024] = 8'h6F;
Memory[21031] = 8'h27;
Memory[21030] = 8'h4D;
Memory[21029] = 8'h21;
Memory[21028] = 8'h83;
Memory[21035] = 8'h00;
Memory[21034] = 8'h3B;
Memory[21033] = 8'h2A;
Memory[21032] = 8'h23;
Memory[21039] = 8'h12;
Memory[21038] = 8'h40;
Memory[21037] = 8'h20;
Memory[21036] = 8'h6F;
Memory[21043] = 8'h27;
Memory[21042] = 8'h8D;
Memory[21041] = 8'h21;
Memory[21040] = 8'h83;
Memory[21047] = 8'h00;
Memory[21046] = 8'h3B;
Memory[21045] = 8'h2A;
Memory[21044] = 8'h23;
Memory[21051] = 8'h12;
Memory[21050] = 8'h40;
Memory[21049] = 8'h20;
Memory[21048] = 8'h6F;
Memory[21055] = 8'h27;
Memory[21054] = 8'hCD;
Memory[21053] = 8'h21;
Memory[21052] = 8'h83;
Memory[21059] = 8'h00;
Memory[21058] = 8'h3B;
Memory[21057] = 8'h2A;
Memory[21056] = 8'h23;
Memory[21063] = 8'h12;
Memory[21062] = 8'h40;
Memory[21061] = 8'h20;
Memory[21060] = 8'h6F;
Memory[21067] = 8'h28;
Memory[21066] = 8'h0D;
Memory[21065] = 8'h21;
Memory[21064] = 8'h83;
Memory[21071] = 8'h00;
Memory[21070] = 8'h3B;
Memory[21069] = 8'h2A;
Memory[21068] = 8'h23;
Memory[21075] = 8'h12;
Memory[21074] = 8'h40;
Memory[21073] = 8'h20;
Memory[21072] = 8'h6F;
Memory[21079] = 8'h28;
Memory[21078] = 8'h4D;
Memory[21077] = 8'h21;
Memory[21076] = 8'h83;
Memory[21083] = 8'h00;
Memory[21082] = 8'h3B;
Memory[21081] = 8'h2A;
Memory[21080] = 8'h23;
Memory[21087] = 8'h12;
Memory[21086] = 8'h40;
Memory[21085] = 8'h20;
Memory[21084] = 8'h6F;
Memory[21091] = 8'h28;
Memory[21090] = 8'h8D;
Memory[21089] = 8'h21;
Memory[21088] = 8'h83;
Memory[21095] = 8'h00;
Memory[21094] = 8'h3B;
Memory[21093] = 8'h2A;
Memory[21092] = 8'h23;
Memory[21099] = 8'h12;
Memory[21098] = 8'h40;
Memory[21097] = 8'h20;
Memory[21096] = 8'h6F;
Memory[21103] = 8'h28;
Memory[21102] = 8'hCD;
Memory[21101] = 8'h21;
Memory[21100] = 8'h83;
Memory[21107] = 8'h00;
Memory[21106] = 8'h3B;
Memory[21105] = 8'h2A;
Memory[21104] = 8'h23;
Memory[21111] = 8'h12;
Memory[21110] = 8'h40;
Memory[21109] = 8'h20;
Memory[21108] = 8'h6F;
Memory[21115] = 8'h29;
Memory[21114] = 8'h0D;
Memory[21113] = 8'h21;
Memory[21112] = 8'h83;
Memory[21119] = 8'h00;
Memory[21118] = 8'h3B;
Memory[21117] = 8'h2A;
Memory[21116] = 8'h23;
Memory[21123] = 8'h12;
Memory[21122] = 8'h40;
Memory[21121] = 8'h20;
Memory[21120] = 8'h6F;
Memory[21127] = 8'h29;
Memory[21126] = 8'h4D;
Memory[21125] = 8'h21;
Memory[21124] = 8'h83;
Memory[21131] = 8'h00;
Memory[21130] = 8'h3B;
Memory[21129] = 8'h2A;
Memory[21128] = 8'h23;
Memory[21135] = 8'h12;
Memory[21134] = 8'h40;
Memory[21133] = 8'h20;
Memory[21132] = 8'h6F;
Memory[21139] = 8'h29;
Memory[21138] = 8'h8D;
Memory[21137] = 8'h21;
Memory[21136] = 8'h83;
Memory[21143] = 8'h00;
Memory[21142] = 8'h3B;
Memory[21141] = 8'h2A;
Memory[21140] = 8'h23;
Memory[21147] = 8'h12;
Memory[21146] = 8'h40;
Memory[21145] = 8'h20;
Memory[21144] = 8'h6F;
Memory[21151] = 8'h29;
Memory[21150] = 8'hCD;
Memory[21149] = 8'h21;
Memory[21148] = 8'h83;
Memory[21155] = 8'h00;
Memory[21154] = 8'h3B;
Memory[21153] = 8'h2A;
Memory[21152] = 8'h23;
Memory[21159] = 8'h12;
Memory[21158] = 8'h40;
Memory[21157] = 8'h20;
Memory[21156] = 8'h6F;
Memory[21163] = 8'h2A;
Memory[21162] = 8'h0D;
Memory[21161] = 8'h21;
Memory[21160] = 8'h83;
Memory[21167] = 8'h00;
Memory[21166] = 8'h3B;
Memory[21165] = 8'h2A;
Memory[21164] = 8'h23;
Memory[21171] = 8'h12;
Memory[21170] = 8'h40;
Memory[21169] = 8'h20;
Memory[21168] = 8'h6F;
Memory[21175] = 8'h2A;
Memory[21174] = 8'h4D;
Memory[21173] = 8'h21;
Memory[21172] = 8'h83;
Memory[21179] = 8'h00;
Memory[21178] = 8'h3B;
Memory[21177] = 8'h2A;
Memory[21176] = 8'h23;
Memory[21183] = 8'h12;
Memory[21182] = 8'h40;
Memory[21181] = 8'h20;
Memory[21180] = 8'h6F;
Memory[21187] = 8'h2A;
Memory[21186] = 8'h8D;
Memory[21185] = 8'h21;
Memory[21184] = 8'h83;
Memory[21191] = 8'h00;
Memory[21190] = 8'h3B;
Memory[21189] = 8'h2A;
Memory[21188] = 8'h23;
Memory[21195] = 8'h12;
Memory[21194] = 8'h40;
Memory[21193] = 8'h20;
Memory[21192] = 8'h6F;
Memory[21199] = 8'h2A;
Memory[21198] = 8'hCD;
Memory[21197] = 8'h21;
Memory[21196] = 8'h83;
Memory[21203] = 8'h00;
Memory[21202] = 8'h3B;
Memory[21201] = 8'h2A;
Memory[21200] = 8'h23;
Memory[21207] = 8'h12;
Memory[21206] = 8'h40;
Memory[21205] = 8'h20;
Memory[21204] = 8'h6F;
Memory[21211] = 8'h2B;
Memory[21210] = 8'h0D;
Memory[21209] = 8'h21;
Memory[21208] = 8'h83;
Memory[21215] = 8'h00;
Memory[21214] = 8'h3B;
Memory[21213] = 8'h2A;
Memory[21212] = 8'h23;
Memory[21219] = 8'h12;
Memory[21218] = 8'h40;
Memory[21217] = 8'h20;
Memory[21216] = 8'h6F;
Memory[21223] = 8'h2B;
Memory[21222] = 8'h4D;
Memory[21221] = 8'h21;
Memory[21220] = 8'h83;
Memory[21227] = 8'h00;
Memory[21226] = 8'h3B;
Memory[21225] = 8'h2A;
Memory[21224] = 8'h23;
Memory[21231] = 8'h12;
Memory[21230] = 8'h40;
Memory[21229] = 8'h20;
Memory[21228] = 8'h6F;
Memory[21235] = 8'h2B;
Memory[21234] = 8'h8D;
Memory[21233] = 8'h21;
Memory[21232] = 8'h83;
Memory[21239] = 8'h00;
Memory[21238] = 8'h3B;
Memory[21237] = 8'h2A;
Memory[21236] = 8'h23;
Memory[21243] = 8'h12;
Memory[21242] = 8'h40;
Memory[21241] = 8'h20;
Memory[21240] = 8'h6F;
Memory[21247] = 8'h2B;
Memory[21246] = 8'hCD;
Memory[21245] = 8'h21;
Memory[21244] = 8'h83;
Memory[21251] = 8'h00;
Memory[21250] = 8'h3B;
Memory[21249] = 8'h2A;
Memory[21248] = 8'h23;
Memory[21255] = 8'h12;
Memory[21254] = 8'h40;
Memory[21253] = 8'h20;
Memory[21252] = 8'h6F;
Memory[21259] = 8'h2C;
Memory[21258] = 8'h0D;
Memory[21257] = 8'h21;
Memory[21256] = 8'h83;
Memory[21263] = 8'h00;
Memory[21262] = 8'h3B;
Memory[21261] = 8'h2A;
Memory[21260] = 8'h23;
Memory[21267] = 8'h12;
Memory[21266] = 8'h40;
Memory[21265] = 8'h20;
Memory[21264] = 8'h6F;
Memory[21271] = 8'h2C;
Memory[21270] = 8'h4D;
Memory[21269] = 8'h21;
Memory[21268] = 8'h83;
Memory[21275] = 8'h00;
Memory[21274] = 8'h3B;
Memory[21273] = 8'h2A;
Memory[21272] = 8'h23;
Memory[21279] = 8'h12;
Memory[21278] = 8'h40;
Memory[21277] = 8'h20;
Memory[21276] = 8'h6F;
Memory[21283] = 8'h2C;
Memory[21282] = 8'h8D;
Memory[21281] = 8'h21;
Memory[21280] = 8'h83;
Memory[21287] = 8'h00;
Memory[21286] = 8'h3B;
Memory[21285] = 8'h2A;
Memory[21284] = 8'h23;
Memory[21291] = 8'h12;
Memory[21290] = 8'h40;
Memory[21289] = 8'h20;
Memory[21288] = 8'h6F;
Memory[21295] = 8'h2C;
Memory[21294] = 8'hCD;
Memory[21293] = 8'h21;
Memory[21292] = 8'h83;
Memory[21299] = 8'h00;
Memory[21298] = 8'h3B;
Memory[21297] = 8'h2A;
Memory[21296] = 8'h23;
Memory[21303] = 8'h12;
Memory[21302] = 8'h40;
Memory[21301] = 8'h20;
Memory[21300] = 8'h6F;
Memory[21307] = 8'h2D;
Memory[21306] = 8'h0D;
Memory[21305] = 8'h21;
Memory[21304] = 8'h83;
Memory[21311] = 8'h00;
Memory[21310] = 8'h3B;
Memory[21309] = 8'h2A;
Memory[21308] = 8'h23;
Memory[21315] = 8'h12;
Memory[21314] = 8'h40;
Memory[21313] = 8'h20;
Memory[21312] = 8'h6F;
Memory[21319] = 8'h2D;
Memory[21318] = 8'h4D;
Memory[21317] = 8'h21;
Memory[21316] = 8'h83;
Memory[21323] = 8'h00;
Memory[21322] = 8'h3B;
Memory[21321] = 8'h2A;
Memory[21320] = 8'h23;
Memory[21327] = 8'h12;
Memory[21326] = 8'h40;
Memory[21325] = 8'h20;
Memory[21324] = 8'h6F;
Memory[21331] = 8'h2D;
Memory[21330] = 8'h8D;
Memory[21329] = 8'h21;
Memory[21328] = 8'h83;
Memory[21335] = 8'h00;
Memory[21334] = 8'h3B;
Memory[21333] = 8'h2A;
Memory[21332] = 8'h23;
Memory[21339] = 8'h12;
Memory[21338] = 8'h40;
Memory[21337] = 8'h20;
Memory[21336] = 8'h6F;
Memory[21343] = 8'h2D;
Memory[21342] = 8'hCD;
Memory[21341] = 8'h21;
Memory[21340] = 8'h83;
Memory[21347] = 8'h00;
Memory[21346] = 8'h3B;
Memory[21345] = 8'h2A;
Memory[21344] = 8'h23;
Memory[21351] = 8'h12;
Memory[21350] = 8'h40;
Memory[21349] = 8'h20;
Memory[21348] = 8'h6F;
Memory[21355] = 8'h2E;
Memory[21354] = 8'h0D;
Memory[21353] = 8'h21;
Memory[21352] = 8'h83;
Memory[21359] = 8'h00;
Memory[21358] = 8'h3B;
Memory[21357] = 8'h2A;
Memory[21356] = 8'h23;
Memory[21363] = 8'h12;
Memory[21362] = 8'h40;
Memory[21361] = 8'h20;
Memory[21360] = 8'h6F;
Memory[21367] = 8'h2E;
Memory[21366] = 8'h4D;
Memory[21365] = 8'h21;
Memory[21364] = 8'h83;
Memory[21371] = 8'h00;
Memory[21370] = 8'h3B;
Memory[21369] = 8'h2A;
Memory[21368] = 8'h23;
Memory[21375] = 8'h12;
Memory[21374] = 8'h40;
Memory[21373] = 8'h20;
Memory[21372] = 8'h6F;
Memory[21379] = 8'h2E;
Memory[21378] = 8'h8D;
Memory[21377] = 8'h21;
Memory[21376] = 8'h83;
Memory[21383] = 8'h00;
Memory[21382] = 8'h3B;
Memory[21381] = 8'h2A;
Memory[21380] = 8'h23;
Memory[21387] = 8'h12;
Memory[21386] = 8'h40;
Memory[21385] = 8'h20;
Memory[21384] = 8'h6F;
Memory[21391] = 8'h2E;
Memory[21390] = 8'hCD;
Memory[21389] = 8'h21;
Memory[21388] = 8'h83;
Memory[21395] = 8'h00;
Memory[21394] = 8'h3B;
Memory[21393] = 8'h2A;
Memory[21392] = 8'h23;
Memory[21399] = 8'h12;
Memory[21398] = 8'h40;
Memory[21397] = 8'h20;
Memory[21396] = 8'h6F;
Memory[21403] = 8'h2F;
Memory[21402] = 8'h0D;
Memory[21401] = 8'h21;
Memory[21400] = 8'h83;
Memory[21407] = 8'h00;
Memory[21406] = 8'h3B;
Memory[21405] = 8'h2A;
Memory[21404] = 8'h23;
Memory[21411] = 8'h12;
Memory[21410] = 8'h40;
Memory[21409] = 8'h20;
Memory[21408] = 8'h6F;
Memory[21415] = 8'h2F;
Memory[21414] = 8'h4D;
Memory[21413] = 8'h21;
Memory[21412] = 8'h83;
Memory[21419] = 8'h00;
Memory[21418] = 8'h3B;
Memory[21417] = 8'h2A;
Memory[21416] = 8'h23;
Memory[21423] = 8'h12;
Memory[21422] = 8'h40;
Memory[21421] = 8'h20;
Memory[21420] = 8'h6F;
Memory[21427] = 8'h2F;
Memory[21426] = 8'h8D;
Memory[21425] = 8'h21;
Memory[21424] = 8'h83;
Memory[21431] = 8'h00;
Memory[21430] = 8'h3B;
Memory[21429] = 8'h2A;
Memory[21428] = 8'h23;
Memory[21435] = 8'h12;
Memory[21434] = 8'h40;
Memory[21433] = 8'h20;
Memory[21432] = 8'h6F;
Memory[21439] = 8'h2F;
Memory[21438] = 8'hCD;
Memory[21437] = 8'h21;
Memory[21436] = 8'h83;
Memory[21443] = 8'h00;
Memory[21442] = 8'h3B;
Memory[21441] = 8'h2A;
Memory[21440] = 8'h23;
Memory[21447] = 8'h12;
Memory[21446] = 8'h40;
Memory[21445] = 8'h20;
Memory[21444] = 8'h6F;
Memory[21451] = 8'h30;
Memory[21450] = 8'h0D;
Memory[21449] = 8'h21;
Memory[21448] = 8'h83;
Memory[21455] = 8'h00;
Memory[21454] = 8'h3B;
Memory[21453] = 8'h2A;
Memory[21452] = 8'h23;
Memory[21459] = 8'h12;
Memory[21458] = 8'h40;
Memory[21457] = 8'h20;
Memory[21456] = 8'h6F;
Memory[21463] = 8'h30;
Memory[21462] = 8'h4D;
Memory[21461] = 8'h21;
Memory[21460] = 8'h83;
Memory[21467] = 8'h00;
Memory[21466] = 8'h3B;
Memory[21465] = 8'h2A;
Memory[21464] = 8'h23;
Memory[21471] = 8'h12;
Memory[21470] = 8'h40;
Memory[21469] = 8'h20;
Memory[21468] = 8'h6F;
Memory[21475] = 8'h30;
Memory[21474] = 8'h8D;
Memory[21473] = 8'h21;
Memory[21472] = 8'h83;
Memory[21479] = 8'h00;
Memory[21478] = 8'h3B;
Memory[21477] = 8'h2A;
Memory[21476] = 8'h23;
Memory[21483] = 8'h12;
Memory[21482] = 8'h40;
Memory[21481] = 8'h20;
Memory[21480] = 8'h6F;
Memory[21487] = 8'h30;
Memory[21486] = 8'hCD;
Memory[21485] = 8'h21;
Memory[21484] = 8'h83;
Memory[21491] = 8'h00;
Memory[21490] = 8'h3B;
Memory[21489] = 8'h2A;
Memory[21488] = 8'h23;
Memory[21495] = 8'h12;
Memory[21494] = 8'h40;
Memory[21493] = 8'h20;
Memory[21492] = 8'h6F;
Memory[21499] = 8'h31;
Memory[21498] = 8'h0D;
Memory[21497] = 8'h21;
Memory[21496] = 8'h83;
Memory[21503] = 8'h00;
Memory[21502] = 8'h3B;
Memory[21501] = 8'h2A;
Memory[21500] = 8'h23;
Memory[21507] = 8'h12;
Memory[21506] = 8'h40;
Memory[21505] = 8'h20;
Memory[21504] = 8'h6F;
Memory[21511] = 8'h31;
Memory[21510] = 8'h4D;
Memory[21509] = 8'h21;
Memory[21508] = 8'h83;
Memory[21515] = 8'h00;
Memory[21514] = 8'h3B;
Memory[21513] = 8'h2A;
Memory[21512] = 8'h23;
Memory[21519] = 8'h12;
Memory[21518] = 8'h40;
Memory[21517] = 8'h20;
Memory[21516] = 8'h6F;
Memory[21523] = 8'h31;
Memory[21522] = 8'h8D;
Memory[21521] = 8'h21;
Memory[21520] = 8'h83;
Memory[21527] = 8'h00;
Memory[21526] = 8'h3B;
Memory[21525] = 8'h2A;
Memory[21524] = 8'h23;
Memory[21531] = 8'h12;
Memory[21530] = 8'h40;
Memory[21529] = 8'h20;
Memory[21528] = 8'h6F;
Memory[21535] = 8'h31;
Memory[21534] = 8'hCD;
Memory[21533] = 8'h21;
Memory[21532] = 8'h83;
Memory[21539] = 8'h00;
Memory[21538] = 8'h3B;
Memory[21537] = 8'h2A;
Memory[21536] = 8'h23;
Memory[21543] = 8'h12;
Memory[21542] = 8'h40;
Memory[21541] = 8'h20;
Memory[21540] = 8'h6F;
Memory[21547] = 8'h32;
Memory[21546] = 8'h0D;
Memory[21545] = 8'h21;
Memory[21544] = 8'h83;
Memory[21551] = 8'h00;
Memory[21550] = 8'h3B;
Memory[21549] = 8'h2A;
Memory[21548] = 8'h23;
Memory[21555] = 8'h12;
Memory[21554] = 8'h40;
Memory[21553] = 8'h20;
Memory[21552] = 8'h6F;
Memory[21559] = 8'h32;
Memory[21558] = 8'h4D;
Memory[21557] = 8'h21;
Memory[21556] = 8'h83;
Memory[21563] = 8'h00;
Memory[21562] = 8'h3B;
Memory[21561] = 8'h2A;
Memory[21560] = 8'h23;
Memory[21567] = 8'h12;
Memory[21566] = 8'h40;
Memory[21565] = 8'h20;
Memory[21564] = 8'h6F;
Memory[21571] = 8'h32;
Memory[21570] = 8'h8D;
Memory[21569] = 8'h21;
Memory[21568] = 8'h83;
Memory[21575] = 8'h00;
Memory[21574] = 8'h3B;
Memory[21573] = 8'h2A;
Memory[21572] = 8'h23;
Memory[21579] = 8'h12;
Memory[21578] = 8'h40;
Memory[21577] = 8'h20;
Memory[21576] = 8'h6F;
Memory[21583] = 8'h32;
Memory[21582] = 8'hCD;
Memory[21581] = 8'h21;
Memory[21580] = 8'h83;
Memory[21587] = 8'h00;
Memory[21586] = 8'h3B;
Memory[21585] = 8'h2A;
Memory[21584] = 8'h23;
Memory[21591] = 8'h12;
Memory[21590] = 8'h40;
Memory[21589] = 8'h20;
Memory[21588] = 8'h6F;
Memory[21595] = 8'h33;
Memory[21594] = 8'h0D;
Memory[21593] = 8'h21;
Memory[21592] = 8'h83;
Memory[21599] = 8'h00;
Memory[21598] = 8'h3B;
Memory[21597] = 8'h2A;
Memory[21596] = 8'h23;
Memory[21603] = 8'h12;
Memory[21602] = 8'h40;
Memory[21601] = 8'h20;
Memory[21600] = 8'h6F;
Memory[21607] = 8'h33;
Memory[21606] = 8'h4D;
Memory[21605] = 8'h21;
Memory[21604] = 8'h83;
Memory[21611] = 8'h00;
Memory[21610] = 8'h3B;
Memory[21609] = 8'h2A;
Memory[21608] = 8'h23;
Memory[21615] = 8'h12;
Memory[21614] = 8'h40;
Memory[21613] = 8'h20;
Memory[21612] = 8'h6F;
Memory[21619] = 8'h33;
Memory[21618] = 8'h8D;
Memory[21617] = 8'h21;
Memory[21616] = 8'h83;
Memory[21623] = 8'h00;
Memory[21622] = 8'h3B;
Memory[21621] = 8'h2A;
Memory[21620] = 8'h23;
Memory[21627] = 8'h12;
Memory[21626] = 8'h40;
Memory[21625] = 8'h20;
Memory[21624] = 8'h6F;
Memory[21631] = 8'h33;
Memory[21630] = 8'hCD;
Memory[21629] = 8'h21;
Memory[21628] = 8'h83;
Memory[21635] = 8'h00;
Memory[21634] = 8'h3B;
Memory[21633] = 8'h2A;
Memory[21632] = 8'h23;
Memory[21639] = 8'h12;
Memory[21638] = 8'h40;
Memory[21637] = 8'h20;
Memory[21636] = 8'h6F;
Memory[21643] = 8'h34;
Memory[21642] = 8'h0D;
Memory[21641] = 8'h21;
Memory[21640] = 8'h83;
Memory[21647] = 8'h00;
Memory[21646] = 8'h3B;
Memory[21645] = 8'h2A;
Memory[21644] = 8'h23;
Memory[21651] = 8'h12;
Memory[21650] = 8'h40;
Memory[21649] = 8'h20;
Memory[21648] = 8'h6F;
Memory[21655] = 8'h34;
Memory[21654] = 8'h4D;
Memory[21653] = 8'h21;
Memory[21652] = 8'h83;
Memory[21659] = 8'h00;
Memory[21658] = 8'h3B;
Memory[21657] = 8'h2A;
Memory[21656] = 8'h23;
Memory[21663] = 8'h12;
Memory[21662] = 8'h40;
Memory[21661] = 8'h20;
Memory[21660] = 8'h6F;
Memory[21667] = 8'h34;
Memory[21666] = 8'h8D;
Memory[21665] = 8'h21;
Memory[21664] = 8'h83;
Memory[21671] = 8'h00;
Memory[21670] = 8'h3B;
Memory[21669] = 8'h2A;
Memory[21668] = 8'h23;
Memory[21675] = 8'h12;
Memory[21674] = 8'h40;
Memory[21673] = 8'h20;
Memory[21672] = 8'h6F;
Memory[21679] = 8'h34;
Memory[21678] = 8'hCD;
Memory[21677] = 8'h21;
Memory[21676] = 8'h83;
Memory[21683] = 8'h00;
Memory[21682] = 8'h3B;
Memory[21681] = 8'h2A;
Memory[21680] = 8'h23;
Memory[21687] = 8'h12;
Memory[21686] = 8'h40;
Memory[21685] = 8'h20;
Memory[21684] = 8'h6F;
Memory[21691] = 8'h35;
Memory[21690] = 8'h0D;
Memory[21689] = 8'h21;
Memory[21688] = 8'h83;
Memory[21695] = 8'h00;
Memory[21694] = 8'h3B;
Memory[21693] = 8'h2A;
Memory[21692] = 8'h23;
Memory[21699] = 8'h12;
Memory[21698] = 8'h40;
Memory[21697] = 8'h20;
Memory[21696] = 8'h6F;
Memory[21703] = 8'h35;
Memory[21702] = 8'h4D;
Memory[21701] = 8'h21;
Memory[21700] = 8'h83;
Memory[21707] = 8'h00;
Memory[21706] = 8'h3B;
Memory[21705] = 8'h2A;
Memory[21704] = 8'h23;
Memory[21711] = 8'h12;
Memory[21710] = 8'h40;
Memory[21709] = 8'h20;
Memory[21708] = 8'h6F;
Memory[21715] = 8'h35;
Memory[21714] = 8'h8D;
Memory[21713] = 8'h21;
Memory[21712] = 8'h83;
Memory[21719] = 8'h00;
Memory[21718] = 8'h3B;
Memory[21717] = 8'h2A;
Memory[21716] = 8'h23;
Memory[21723] = 8'h12;
Memory[21722] = 8'h40;
Memory[21721] = 8'h20;
Memory[21720] = 8'h6F;
Memory[21727] = 8'h35;
Memory[21726] = 8'hCD;
Memory[21725] = 8'h21;
Memory[21724] = 8'h83;
Memory[21731] = 8'h00;
Memory[21730] = 8'h3B;
Memory[21729] = 8'h2A;
Memory[21728] = 8'h23;
Memory[21735] = 8'h12;
Memory[21734] = 8'h40;
Memory[21733] = 8'h20;
Memory[21732] = 8'h6F;
Memory[21739] = 8'h36;
Memory[21738] = 8'h0D;
Memory[21737] = 8'h21;
Memory[21736] = 8'h83;
Memory[21743] = 8'h00;
Memory[21742] = 8'h3B;
Memory[21741] = 8'h2A;
Memory[21740] = 8'h23;
Memory[21747] = 8'h12;
Memory[21746] = 8'h40;
Memory[21745] = 8'h20;
Memory[21744] = 8'h6F;
Memory[21751] = 8'h36;
Memory[21750] = 8'h4D;
Memory[21749] = 8'h21;
Memory[21748] = 8'h83;
Memory[21755] = 8'h00;
Memory[21754] = 8'h3B;
Memory[21753] = 8'h2A;
Memory[21752] = 8'h23;
Memory[21759] = 8'h12;
Memory[21758] = 8'h40;
Memory[21757] = 8'h20;
Memory[21756] = 8'h6F;
Memory[21763] = 8'h36;
Memory[21762] = 8'h8D;
Memory[21761] = 8'h21;
Memory[21760] = 8'h83;
Memory[21767] = 8'h00;
Memory[21766] = 8'h3B;
Memory[21765] = 8'h2A;
Memory[21764] = 8'h23;
Memory[21771] = 8'h12;
Memory[21770] = 8'h40;
Memory[21769] = 8'h20;
Memory[21768] = 8'h6F;
Memory[21775] = 8'h36;
Memory[21774] = 8'hCD;
Memory[21773] = 8'h21;
Memory[21772] = 8'h83;
Memory[21779] = 8'h00;
Memory[21778] = 8'h3B;
Memory[21777] = 8'h2A;
Memory[21776] = 8'h23;
Memory[21783] = 8'h12;
Memory[21782] = 8'h40;
Memory[21781] = 8'h20;
Memory[21780] = 8'h6F;
Memory[21787] = 8'h37;
Memory[21786] = 8'h0D;
Memory[21785] = 8'h21;
Memory[21784] = 8'h83;
Memory[21791] = 8'h00;
Memory[21790] = 8'h3B;
Memory[21789] = 8'h2A;
Memory[21788] = 8'h23;
Memory[21795] = 8'h12;
Memory[21794] = 8'h40;
Memory[21793] = 8'h20;
Memory[21792] = 8'h6F;
Memory[21799] = 8'h37;
Memory[21798] = 8'h4D;
Memory[21797] = 8'h21;
Memory[21796] = 8'h83;
Memory[21803] = 8'h00;
Memory[21802] = 8'h3B;
Memory[21801] = 8'h2A;
Memory[21800] = 8'h23;
Memory[21807] = 8'h12;
Memory[21806] = 8'h40;
Memory[21805] = 8'h20;
Memory[21804] = 8'h6F;
Memory[21811] = 8'h37;
Memory[21810] = 8'h8D;
Memory[21809] = 8'h21;
Memory[21808] = 8'h83;
Memory[21815] = 8'h00;
Memory[21814] = 8'h3B;
Memory[21813] = 8'h2A;
Memory[21812] = 8'h23;
Memory[21819] = 8'h12;
Memory[21818] = 8'h40;
Memory[21817] = 8'h20;
Memory[21816] = 8'h6F;
Memory[21823] = 8'h37;
Memory[21822] = 8'hCD;
Memory[21821] = 8'h21;
Memory[21820] = 8'h83;
Memory[21827] = 8'h00;
Memory[21826] = 8'h3B;
Memory[21825] = 8'h2A;
Memory[21824] = 8'h23;
Memory[21831] = 8'h12;
Memory[21830] = 8'h40;
Memory[21829] = 8'h20;
Memory[21828] = 8'h6F;
Memory[21835] = 8'h38;
Memory[21834] = 8'h0D;
Memory[21833] = 8'h21;
Memory[21832] = 8'h83;
Memory[21839] = 8'h00;
Memory[21838] = 8'h3B;
Memory[21837] = 8'h2A;
Memory[21836] = 8'h23;
Memory[21843] = 8'h12;
Memory[21842] = 8'h40;
Memory[21841] = 8'h20;
Memory[21840] = 8'h6F;
Memory[21847] = 8'h38;
Memory[21846] = 8'h4D;
Memory[21845] = 8'h21;
Memory[21844] = 8'h83;
Memory[21851] = 8'h00;
Memory[21850] = 8'h3B;
Memory[21849] = 8'h2A;
Memory[21848] = 8'h23;
Memory[21855] = 8'h12;
Memory[21854] = 8'h40;
Memory[21853] = 8'h20;
Memory[21852] = 8'h6F;
Memory[21859] = 8'h38;
Memory[21858] = 8'h8D;
Memory[21857] = 8'h21;
Memory[21856] = 8'h83;
Memory[21863] = 8'h00;
Memory[21862] = 8'h3B;
Memory[21861] = 8'h2A;
Memory[21860] = 8'h23;
Memory[21867] = 8'h12;
Memory[21866] = 8'h40;
Memory[21865] = 8'h20;
Memory[21864] = 8'h6F;
Memory[21871] = 8'h38;
Memory[21870] = 8'hCD;
Memory[21869] = 8'h21;
Memory[21868] = 8'h83;
Memory[21875] = 8'h00;
Memory[21874] = 8'h3B;
Memory[21873] = 8'h2A;
Memory[21872] = 8'h23;
Memory[21879] = 8'h12;
Memory[21878] = 8'h40;
Memory[21877] = 8'h20;
Memory[21876] = 8'h6F;
Memory[21883] = 8'h39;
Memory[21882] = 8'h0D;
Memory[21881] = 8'h21;
Memory[21880] = 8'h83;
Memory[21887] = 8'h00;
Memory[21886] = 8'h3B;
Memory[21885] = 8'h2A;
Memory[21884] = 8'h23;
Memory[21891] = 8'h12;
Memory[21890] = 8'h40;
Memory[21889] = 8'h20;
Memory[21888] = 8'h6F;
Memory[21895] = 8'h39;
Memory[21894] = 8'h4D;
Memory[21893] = 8'h21;
Memory[21892] = 8'h83;
Memory[21899] = 8'h00;
Memory[21898] = 8'h3B;
Memory[21897] = 8'h2A;
Memory[21896] = 8'h23;
Memory[21903] = 8'h12;
Memory[21902] = 8'h40;
Memory[21901] = 8'h20;
Memory[21900] = 8'h6F;
Memory[21907] = 8'h39;
Memory[21906] = 8'h8D;
Memory[21905] = 8'h21;
Memory[21904] = 8'h83;
Memory[21911] = 8'h00;
Memory[21910] = 8'h3B;
Memory[21909] = 8'h2A;
Memory[21908] = 8'h23;
Memory[21915] = 8'h12;
Memory[21914] = 8'h40;
Memory[21913] = 8'h20;
Memory[21912] = 8'h6F;
Memory[21919] = 8'h39;
Memory[21918] = 8'hCD;
Memory[21917] = 8'h21;
Memory[21916] = 8'h83;
Memory[21923] = 8'h00;
Memory[21922] = 8'h3B;
Memory[21921] = 8'h2A;
Memory[21920] = 8'h23;
Memory[21927] = 8'h12;
Memory[21926] = 8'h40;
Memory[21925] = 8'h20;
Memory[21924] = 8'h6F;
Memory[21931] = 8'h3A;
Memory[21930] = 8'h0D;
Memory[21929] = 8'h21;
Memory[21928] = 8'h83;
Memory[21935] = 8'h00;
Memory[21934] = 8'h3B;
Memory[21933] = 8'h2A;
Memory[21932] = 8'h23;
Memory[21939] = 8'h12;
Memory[21938] = 8'h40;
Memory[21937] = 8'h20;
Memory[21936] = 8'h6F;
Memory[21943] = 8'h3A;
Memory[21942] = 8'h4D;
Memory[21941] = 8'h21;
Memory[21940] = 8'h83;
Memory[21947] = 8'h00;
Memory[21946] = 8'h3B;
Memory[21945] = 8'h2A;
Memory[21944] = 8'h23;
Memory[21951] = 8'h12;
Memory[21950] = 8'h40;
Memory[21949] = 8'h20;
Memory[21948] = 8'h6F;
Memory[21955] = 8'h3A;
Memory[21954] = 8'h8D;
Memory[21953] = 8'h21;
Memory[21952] = 8'h83;
Memory[21959] = 8'h00;
Memory[21958] = 8'h3B;
Memory[21957] = 8'h2A;
Memory[21956] = 8'h23;
Memory[21963] = 8'h12;
Memory[21962] = 8'h40;
Memory[21961] = 8'h20;
Memory[21960] = 8'h6F;
Memory[21967] = 8'h3A;
Memory[21966] = 8'hCD;
Memory[21965] = 8'h21;
Memory[21964] = 8'h83;
Memory[21971] = 8'h00;
Memory[21970] = 8'h3B;
Memory[21969] = 8'h2A;
Memory[21968] = 8'h23;
Memory[21975] = 8'h12;
Memory[21974] = 8'h40;
Memory[21973] = 8'h20;
Memory[21972] = 8'h6F;
Memory[21979] = 8'h3B;
Memory[21978] = 8'h0D;
Memory[21977] = 8'h21;
Memory[21976] = 8'h83;
Memory[21983] = 8'h00;
Memory[21982] = 8'h3B;
Memory[21981] = 8'h2A;
Memory[21980] = 8'h23;
Memory[21987] = 8'h12;
Memory[21986] = 8'h40;
Memory[21985] = 8'h20;
Memory[21984] = 8'h6F;
Memory[21991] = 8'h3B;
Memory[21990] = 8'h4D;
Memory[21989] = 8'h21;
Memory[21988] = 8'h83;
Memory[21995] = 8'h00;
Memory[21994] = 8'h3B;
Memory[21993] = 8'h2A;
Memory[21992] = 8'h23;
Memory[21999] = 8'h12;
Memory[21998] = 8'h40;
Memory[21997] = 8'h20;
Memory[21996] = 8'h6F;
Memory[22003] = 8'h3B;
Memory[22002] = 8'h8D;
Memory[22001] = 8'h21;
Memory[22000] = 8'h83;
Memory[22007] = 8'h00;
Memory[22006] = 8'h3B;
Memory[22005] = 8'h2A;
Memory[22004] = 8'h23;
Memory[22011] = 8'h12;
Memory[22010] = 8'h40;
Memory[22009] = 8'h20;
Memory[22008] = 8'h6F;
Memory[22015] = 8'h3B;
Memory[22014] = 8'hCD;
Memory[22013] = 8'h21;
Memory[22012] = 8'h83;
Memory[22019] = 8'h00;
Memory[22018] = 8'h3B;
Memory[22017] = 8'h2A;
Memory[22016] = 8'h23;
Memory[22023] = 8'h12;
Memory[22022] = 8'h40;
Memory[22021] = 8'h20;
Memory[22020] = 8'h6F;
Memory[22027] = 8'h3C;
Memory[22026] = 8'h0D;
Memory[22025] = 8'h21;
Memory[22024] = 8'h83;
Memory[22031] = 8'h00;
Memory[22030] = 8'h3B;
Memory[22029] = 8'h2A;
Memory[22028] = 8'h23;
Memory[22035] = 8'h12;
Memory[22034] = 8'h40;
Memory[22033] = 8'h20;
Memory[22032] = 8'h6F;
Memory[22039] = 8'h3C;
Memory[22038] = 8'h4D;
Memory[22037] = 8'h21;
Memory[22036] = 8'h83;
Memory[22043] = 8'h00;
Memory[22042] = 8'h3B;
Memory[22041] = 8'h2A;
Memory[22040] = 8'h23;
Memory[22047] = 8'h12;
Memory[22046] = 8'h40;
Memory[22045] = 8'h20;
Memory[22044] = 8'h6F;
Memory[22051] = 8'h3C;
Memory[22050] = 8'h8D;
Memory[22049] = 8'h21;
Memory[22048] = 8'h83;
Memory[22055] = 8'h00;
Memory[22054] = 8'h3B;
Memory[22053] = 8'h2A;
Memory[22052] = 8'h23;
Memory[22059] = 8'h12;
Memory[22058] = 8'h40;
Memory[22057] = 8'h20;
Memory[22056] = 8'h6F;
Memory[22063] = 8'h3C;
Memory[22062] = 8'hCD;
Memory[22061] = 8'h21;
Memory[22060] = 8'h83;
Memory[22067] = 8'h00;
Memory[22066] = 8'h3B;
Memory[22065] = 8'h2A;
Memory[22064] = 8'h23;
Memory[22071] = 8'h12;
Memory[22070] = 8'h40;
Memory[22069] = 8'h20;
Memory[22068] = 8'h6F;
Memory[22075] = 8'h3D;
Memory[22074] = 8'h0D;
Memory[22073] = 8'h21;
Memory[22072] = 8'h83;
Memory[22079] = 8'h00;
Memory[22078] = 8'h3B;
Memory[22077] = 8'h2A;
Memory[22076] = 8'h23;
Memory[22083] = 8'h12;
Memory[22082] = 8'h40;
Memory[22081] = 8'h20;
Memory[22080] = 8'h6F;
Memory[22087] = 8'h3D;
Memory[22086] = 8'h4D;
Memory[22085] = 8'h21;
Memory[22084] = 8'h83;
Memory[22091] = 8'h00;
Memory[22090] = 8'h3B;
Memory[22089] = 8'h2A;
Memory[22088] = 8'h23;
Memory[22095] = 8'h12;
Memory[22094] = 8'h40;
Memory[22093] = 8'h20;
Memory[22092] = 8'h6F;
Memory[22099] = 8'h3D;
Memory[22098] = 8'h8D;
Memory[22097] = 8'h21;
Memory[22096] = 8'h83;
Memory[22103] = 8'h00;
Memory[22102] = 8'h3B;
Memory[22101] = 8'h2A;
Memory[22100] = 8'h23;
Memory[22107] = 8'h12;
Memory[22106] = 8'h40;
Memory[22105] = 8'h20;
Memory[22104] = 8'h6F;
Memory[22111] = 8'h3D;
Memory[22110] = 8'hCD;
Memory[22109] = 8'h21;
Memory[22108] = 8'h83;
Memory[22115] = 8'h00;
Memory[22114] = 8'h3B;
Memory[22113] = 8'h2A;
Memory[22112] = 8'h23;
Memory[22119] = 8'h12;
Memory[22118] = 8'h40;
Memory[22117] = 8'h20;
Memory[22116] = 8'h6F;
Memory[22123] = 8'h3E;
Memory[22122] = 8'h0D;
Memory[22121] = 8'h21;
Memory[22120] = 8'h83;
Memory[22127] = 8'h00;
Memory[22126] = 8'h3B;
Memory[22125] = 8'h2A;
Memory[22124] = 8'h23;
Memory[22131] = 8'h12;
Memory[22130] = 8'h40;
Memory[22129] = 8'h20;
Memory[22128] = 8'h6F;
Memory[22135] = 8'h3E;
Memory[22134] = 8'h4D;
Memory[22133] = 8'h21;
Memory[22132] = 8'h83;
Memory[22139] = 8'h00;
Memory[22138] = 8'h3B;
Memory[22137] = 8'h2A;
Memory[22136] = 8'h23;
Memory[22143] = 8'h12;
Memory[22142] = 8'h40;
Memory[22141] = 8'h20;
Memory[22140] = 8'h6F;
Memory[22147] = 8'h3E;
Memory[22146] = 8'h8D;
Memory[22145] = 8'h21;
Memory[22144] = 8'h83;
Memory[22151] = 8'h00;
Memory[22150] = 8'h3B;
Memory[22149] = 8'h2A;
Memory[22148] = 8'h23;
Memory[22155] = 8'h12;
Memory[22154] = 8'h40;
Memory[22153] = 8'h20;
Memory[22152] = 8'h6F;
Memory[22159] = 8'h3E;
Memory[22158] = 8'hCD;
Memory[22157] = 8'h21;
Memory[22156] = 8'h83;
Memory[22163] = 8'h00;
Memory[22162] = 8'h3B;
Memory[22161] = 8'h2A;
Memory[22160] = 8'h23;
Memory[22167] = 8'h12;
Memory[22166] = 8'h40;
Memory[22165] = 8'h20;
Memory[22164] = 8'h6F;
Memory[22171] = 8'h3F;
Memory[22170] = 8'h0D;
Memory[22169] = 8'h21;
Memory[22168] = 8'h83;
Memory[22175] = 8'h00;
Memory[22174] = 8'h3B;
Memory[22173] = 8'h2A;
Memory[22172] = 8'h23;
Memory[22179] = 8'h12;
Memory[22178] = 8'h40;
Memory[22177] = 8'h20;
Memory[22176] = 8'h6F;
Memory[22183] = 8'h3F;
Memory[22182] = 8'h4D;
Memory[22181] = 8'h21;
Memory[22180] = 8'h83;
Memory[22187] = 8'h00;
Memory[22186] = 8'h3B;
Memory[22185] = 8'h2A;
Memory[22184] = 8'h23;
Memory[22191] = 8'h12;
Memory[22190] = 8'h40;
Memory[22189] = 8'h20;
Memory[22188] = 8'h6F;
Memory[22195] = 8'h3F;
Memory[22194] = 8'h8D;
Memory[22193] = 8'h21;
Memory[22192] = 8'h83;
Memory[22199] = 8'h00;
Memory[22198] = 8'h3B;
Memory[22197] = 8'h2A;
Memory[22196] = 8'h23;
Memory[22203] = 8'h12;
Memory[22202] = 8'h40;
Memory[22201] = 8'h20;
Memory[22200] = 8'h6F;
Memory[22207] = 8'h3F;
Memory[22206] = 8'hCD;
Memory[22205] = 8'h21;
Memory[22204] = 8'h83;
Memory[22211] = 8'h00;
Memory[22210] = 8'h3B;
Memory[22209] = 8'h2A;
Memory[22208] = 8'h23;
Memory[22215] = 8'h12;
Memory[22214] = 8'h40;
Memory[22213] = 8'h20;
Memory[22212] = 8'h6F;
Memory[22219] = 8'h40;
Memory[22218] = 8'h0D;
Memory[22217] = 8'h21;
Memory[22216] = 8'h83;
Memory[22223] = 8'h00;
Memory[22222] = 8'h3B;
Memory[22221] = 8'h2A;
Memory[22220] = 8'h23;
Memory[22227] = 8'h12;
Memory[22226] = 8'h40;
Memory[22225] = 8'h20;
Memory[22224] = 8'h6F;
Memory[22231] = 8'h40;
Memory[22230] = 8'h4D;
Memory[22229] = 8'h21;
Memory[22228] = 8'h83;
Memory[22235] = 8'h00;
Memory[22234] = 8'h3B;
Memory[22233] = 8'h2A;
Memory[22232] = 8'h23;
Memory[22239] = 8'h12;
Memory[22238] = 8'h40;
Memory[22237] = 8'h20;
Memory[22236] = 8'h6F;
Memory[22243] = 8'h40;
Memory[22242] = 8'h8D;
Memory[22241] = 8'h21;
Memory[22240] = 8'h83;
Memory[22247] = 8'h00;
Memory[22246] = 8'h3B;
Memory[22245] = 8'h2A;
Memory[22244] = 8'h23;
Memory[22251] = 8'h12;
Memory[22250] = 8'h40;
Memory[22249] = 8'h20;
Memory[22248] = 8'h6F;
Memory[22255] = 8'h40;
Memory[22254] = 8'hCD;
Memory[22253] = 8'h21;
Memory[22252] = 8'h83;
Memory[22259] = 8'h00;
Memory[22258] = 8'h3B;
Memory[22257] = 8'h2A;
Memory[22256] = 8'h23;
Memory[22263] = 8'h12;
Memory[22262] = 8'h40;
Memory[22261] = 8'h20;
Memory[22260] = 8'h6F;
Memory[22267] = 8'h41;
Memory[22266] = 8'h0D;
Memory[22265] = 8'h21;
Memory[22264] = 8'h83;
Memory[22271] = 8'h00;
Memory[22270] = 8'h3B;
Memory[22269] = 8'h2A;
Memory[22268] = 8'h23;
Memory[22275] = 8'h12;
Memory[22274] = 8'h40;
Memory[22273] = 8'h20;
Memory[22272] = 8'h6F;
Memory[22279] = 8'h41;
Memory[22278] = 8'h4D;
Memory[22277] = 8'h21;
Memory[22276] = 8'h83;
Memory[22283] = 8'h00;
Memory[22282] = 8'h3B;
Memory[22281] = 8'h2A;
Memory[22280] = 8'h23;
Memory[22287] = 8'h12;
Memory[22286] = 8'h40;
Memory[22285] = 8'h20;
Memory[22284] = 8'h6F;
Memory[22291] = 8'h41;
Memory[22290] = 8'h8D;
Memory[22289] = 8'h21;
Memory[22288] = 8'h83;
Memory[22295] = 8'h00;
Memory[22294] = 8'h3B;
Memory[22293] = 8'h2A;
Memory[22292] = 8'h23;
Memory[22299] = 8'h12;
Memory[22298] = 8'h40;
Memory[22297] = 8'h20;
Memory[22296] = 8'h6F;
Memory[22303] = 8'h41;
Memory[22302] = 8'hCD;
Memory[22301] = 8'h21;
Memory[22300] = 8'h83;
Memory[22307] = 8'h00;
Memory[22306] = 8'h3B;
Memory[22305] = 8'h2A;
Memory[22304] = 8'h23;
Memory[22311] = 8'h12;
Memory[22310] = 8'h40;
Memory[22309] = 8'h20;
Memory[22308] = 8'h6F;
Memory[22315] = 8'h42;
Memory[22314] = 8'h0D;
Memory[22313] = 8'h21;
Memory[22312] = 8'h83;
Memory[22319] = 8'h00;
Memory[22318] = 8'h3B;
Memory[22317] = 8'h2A;
Memory[22316] = 8'h23;
Memory[22323] = 8'h12;
Memory[22322] = 8'h40;
Memory[22321] = 8'h20;
Memory[22320] = 8'h6F;
Memory[22327] = 8'h42;
Memory[22326] = 8'h4D;
Memory[22325] = 8'h21;
Memory[22324] = 8'h83;
Memory[22331] = 8'h00;
Memory[22330] = 8'h3B;
Memory[22329] = 8'h2A;
Memory[22328] = 8'h23;
Memory[22335] = 8'h12;
Memory[22334] = 8'h40;
Memory[22333] = 8'h20;
Memory[22332] = 8'h6F;
Memory[22339] = 8'h42;
Memory[22338] = 8'h8D;
Memory[22337] = 8'h21;
Memory[22336] = 8'h83;
Memory[22343] = 8'h00;
Memory[22342] = 8'h3B;
Memory[22341] = 8'h2A;
Memory[22340] = 8'h23;
Memory[22347] = 8'h12;
Memory[22346] = 8'h40;
Memory[22345] = 8'h20;
Memory[22344] = 8'h6F;
Memory[22351] = 8'h42;
Memory[22350] = 8'hCD;
Memory[22349] = 8'h21;
Memory[22348] = 8'h83;
Memory[22355] = 8'h00;
Memory[22354] = 8'h3B;
Memory[22353] = 8'h2A;
Memory[22352] = 8'h23;
Memory[22359] = 8'h12;
Memory[22358] = 8'h40;
Memory[22357] = 8'h20;
Memory[22356] = 8'h6F;
Memory[22363] = 8'h43;
Memory[22362] = 8'h0D;
Memory[22361] = 8'h21;
Memory[22360] = 8'h83;
Memory[22367] = 8'h00;
Memory[22366] = 8'h3B;
Memory[22365] = 8'h2A;
Memory[22364] = 8'h23;
Memory[22371] = 8'h12;
Memory[22370] = 8'h40;
Memory[22369] = 8'h20;
Memory[22368] = 8'h6F;
Memory[22375] = 8'h43;
Memory[22374] = 8'h4D;
Memory[22373] = 8'h21;
Memory[22372] = 8'h83;
Memory[22379] = 8'h00;
Memory[22378] = 8'h3B;
Memory[22377] = 8'h2A;
Memory[22376] = 8'h23;
Memory[22383] = 8'h12;
Memory[22382] = 8'h40;
Memory[22381] = 8'h20;
Memory[22380] = 8'h6F;
Memory[22387] = 8'h43;
Memory[22386] = 8'h8D;
Memory[22385] = 8'h21;
Memory[22384] = 8'h83;
Memory[22391] = 8'h00;
Memory[22390] = 8'h3B;
Memory[22389] = 8'h2A;
Memory[22388] = 8'h23;
Memory[22395] = 8'h12;
Memory[22394] = 8'h40;
Memory[22393] = 8'h20;
Memory[22392] = 8'h6F;
Memory[22399] = 8'h43;
Memory[22398] = 8'hCD;
Memory[22397] = 8'h21;
Memory[22396] = 8'h83;
Memory[22403] = 8'h00;
Memory[22402] = 8'h3B;
Memory[22401] = 8'h2A;
Memory[22400] = 8'h23;
Memory[22407] = 8'h12;
Memory[22406] = 8'h40;
Memory[22405] = 8'h20;
Memory[22404] = 8'h6F;
Memory[22411] = 8'h44;
Memory[22410] = 8'h0D;
Memory[22409] = 8'h21;
Memory[22408] = 8'h83;
Memory[22415] = 8'h00;
Memory[22414] = 8'h3B;
Memory[22413] = 8'h2A;
Memory[22412] = 8'h23;
Memory[22419] = 8'h12;
Memory[22418] = 8'h40;
Memory[22417] = 8'h20;
Memory[22416] = 8'h6F;
Memory[22423] = 8'h44;
Memory[22422] = 8'h4D;
Memory[22421] = 8'h21;
Memory[22420] = 8'h83;
Memory[22427] = 8'h00;
Memory[22426] = 8'h3B;
Memory[22425] = 8'h2A;
Memory[22424] = 8'h23;
Memory[22431] = 8'h12;
Memory[22430] = 8'h40;
Memory[22429] = 8'h20;
Memory[22428] = 8'h6F;
Memory[22435] = 8'h44;
Memory[22434] = 8'h8D;
Memory[22433] = 8'h21;
Memory[22432] = 8'h83;
Memory[22439] = 8'h00;
Memory[22438] = 8'h3B;
Memory[22437] = 8'h2A;
Memory[22436] = 8'h23;
Memory[22443] = 8'h12;
Memory[22442] = 8'h40;
Memory[22441] = 8'h20;
Memory[22440] = 8'h6F;
Memory[22447] = 8'h44;
Memory[22446] = 8'hCD;
Memory[22445] = 8'h21;
Memory[22444] = 8'h83;
Memory[22451] = 8'h00;
Memory[22450] = 8'h3B;
Memory[22449] = 8'h2A;
Memory[22448] = 8'h23;
Memory[22455] = 8'h12;
Memory[22454] = 8'h40;
Memory[22453] = 8'h20;
Memory[22452] = 8'h6F;
Memory[22459] = 8'h45;
Memory[22458] = 8'h0D;
Memory[22457] = 8'h21;
Memory[22456] = 8'h83;
Memory[22463] = 8'h00;
Memory[22462] = 8'h3B;
Memory[22461] = 8'h2A;
Memory[22460] = 8'h23;
Memory[22467] = 8'h12;
Memory[22466] = 8'h40;
Memory[22465] = 8'h20;
Memory[22464] = 8'h6F;
Memory[22471] = 8'h45;
Memory[22470] = 8'h4D;
Memory[22469] = 8'h21;
Memory[22468] = 8'h83;
Memory[22475] = 8'h00;
Memory[22474] = 8'h3B;
Memory[22473] = 8'h2A;
Memory[22472] = 8'h23;
Memory[22479] = 8'h12;
Memory[22478] = 8'h40;
Memory[22477] = 8'h20;
Memory[22476] = 8'h6F;
Memory[22483] = 8'h45;
Memory[22482] = 8'h8D;
Memory[22481] = 8'h21;
Memory[22480] = 8'h83;
Memory[22487] = 8'h00;
Memory[22486] = 8'h3B;
Memory[22485] = 8'h2A;
Memory[22484] = 8'h23;
Memory[22491] = 8'h12;
Memory[22490] = 8'h40;
Memory[22489] = 8'h20;
Memory[22488] = 8'h6F;
Memory[22495] = 8'h45;
Memory[22494] = 8'hCD;
Memory[22493] = 8'h21;
Memory[22492] = 8'h83;
Memory[22499] = 8'h00;
Memory[22498] = 8'h3B;
Memory[22497] = 8'h2A;
Memory[22496] = 8'h23;
Memory[22503] = 8'h12;
Memory[22502] = 8'h40;
Memory[22501] = 8'h20;
Memory[22500] = 8'h6F;
Memory[22507] = 8'h46;
Memory[22506] = 8'h0D;
Memory[22505] = 8'h21;
Memory[22504] = 8'h83;
Memory[22511] = 8'h00;
Memory[22510] = 8'h3B;
Memory[22509] = 8'h2A;
Memory[22508] = 8'h23;
Memory[22515] = 8'h12;
Memory[22514] = 8'h40;
Memory[22513] = 8'h20;
Memory[22512] = 8'h6F;
Memory[22519] = 8'h46;
Memory[22518] = 8'h4D;
Memory[22517] = 8'h21;
Memory[22516] = 8'h83;
Memory[22523] = 8'h00;
Memory[22522] = 8'h3B;
Memory[22521] = 8'h2A;
Memory[22520] = 8'h23;
Memory[22527] = 8'h12;
Memory[22526] = 8'h40;
Memory[22525] = 8'h20;
Memory[22524] = 8'h6F;
Memory[22531] = 8'h46;
Memory[22530] = 8'h8D;
Memory[22529] = 8'h21;
Memory[22528] = 8'h83;
Memory[22535] = 8'h00;
Memory[22534] = 8'h3B;
Memory[22533] = 8'h2A;
Memory[22532] = 8'h23;
Memory[22539] = 8'h12;
Memory[22538] = 8'h40;
Memory[22537] = 8'h20;
Memory[22536] = 8'h6F;
Memory[22543] = 8'h46;
Memory[22542] = 8'hCD;
Memory[22541] = 8'h21;
Memory[22540] = 8'h83;
Memory[22547] = 8'h00;
Memory[22546] = 8'h3B;
Memory[22545] = 8'h2A;
Memory[22544] = 8'h23;
Memory[22551] = 8'h12;
Memory[22550] = 8'h40;
Memory[22549] = 8'h20;
Memory[22548] = 8'h6F;
Memory[22555] = 8'h47;
Memory[22554] = 8'h0D;
Memory[22553] = 8'h21;
Memory[22552] = 8'h83;
Memory[22559] = 8'h00;
Memory[22558] = 8'h3B;
Memory[22557] = 8'h2A;
Memory[22556] = 8'h23;
Memory[22563] = 8'h12;
Memory[22562] = 8'h40;
Memory[22561] = 8'h20;
Memory[22560] = 8'h6F;
Memory[22567] = 8'h47;
Memory[22566] = 8'h4D;
Memory[22565] = 8'h21;
Memory[22564] = 8'h83;
Memory[22571] = 8'h00;
Memory[22570] = 8'h3B;
Memory[22569] = 8'h2A;
Memory[22568] = 8'h23;
Memory[22575] = 8'h12;
Memory[22574] = 8'h40;
Memory[22573] = 8'h20;
Memory[22572] = 8'h6F;
Memory[22579] = 8'h47;
Memory[22578] = 8'h8D;
Memory[22577] = 8'h21;
Memory[22576] = 8'h83;
Memory[22583] = 8'h00;
Memory[22582] = 8'h3B;
Memory[22581] = 8'h2A;
Memory[22580] = 8'h23;
Memory[22587] = 8'h12;
Memory[22586] = 8'h40;
Memory[22585] = 8'h20;
Memory[22584] = 8'h6F;
Memory[22591] = 8'h47;
Memory[22590] = 8'hCD;
Memory[22589] = 8'h21;
Memory[22588] = 8'h83;
Memory[22595] = 8'h00;
Memory[22594] = 8'h3B;
Memory[22593] = 8'h2A;
Memory[22592] = 8'h23;
Memory[22599] = 8'h12;
Memory[22598] = 8'h40;
Memory[22597] = 8'h20;
Memory[22596] = 8'h6F;
Memory[22603] = 8'h48;
Memory[22602] = 8'h0D;
Memory[22601] = 8'h21;
Memory[22600] = 8'h83;
Memory[22607] = 8'h00;
Memory[22606] = 8'h3B;
Memory[22605] = 8'h2A;
Memory[22604] = 8'h23;
Memory[22611] = 8'h12;
Memory[22610] = 8'h40;
Memory[22609] = 8'h20;
Memory[22608] = 8'h6F;
Memory[22615] = 8'h48;
Memory[22614] = 8'h4D;
Memory[22613] = 8'h21;
Memory[22612] = 8'h83;
Memory[22619] = 8'h00;
Memory[22618] = 8'h3B;
Memory[22617] = 8'h2A;
Memory[22616] = 8'h23;
Memory[22623] = 8'h12;
Memory[22622] = 8'h40;
Memory[22621] = 8'h20;
Memory[22620] = 8'h6F;
Memory[22627] = 8'h48;
Memory[22626] = 8'h8D;
Memory[22625] = 8'h21;
Memory[22624] = 8'h83;
Memory[22631] = 8'h00;
Memory[22630] = 8'h3B;
Memory[22629] = 8'h2A;
Memory[22628] = 8'h23;
Memory[22635] = 8'h12;
Memory[22634] = 8'h40;
Memory[22633] = 8'h20;
Memory[22632] = 8'h6F;
Memory[22639] = 8'h48;
Memory[22638] = 8'hCD;
Memory[22637] = 8'h21;
Memory[22636] = 8'h83;
Memory[22643] = 8'h00;
Memory[22642] = 8'h3B;
Memory[22641] = 8'h2A;
Memory[22640] = 8'h23;
Memory[22647] = 8'h12;
Memory[22646] = 8'h40;
Memory[22645] = 8'h20;
Memory[22644] = 8'h6F;
Memory[22651] = 8'h49;
Memory[22650] = 8'h0D;
Memory[22649] = 8'h21;
Memory[22648] = 8'h83;
Memory[22655] = 8'h00;
Memory[22654] = 8'h3B;
Memory[22653] = 8'h2A;
Memory[22652] = 8'h23;
Memory[22659] = 8'h12;
Memory[22658] = 8'h40;
Memory[22657] = 8'h20;
Memory[22656] = 8'h6F;
Memory[22663] = 8'h49;
Memory[22662] = 8'h4D;
Memory[22661] = 8'h21;
Memory[22660] = 8'h83;
Memory[22667] = 8'h00;
Memory[22666] = 8'h3B;
Memory[22665] = 8'h2A;
Memory[22664] = 8'h23;
Memory[22671] = 8'h12;
Memory[22670] = 8'h40;
Memory[22669] = 8'h20;
Memory[22668] = 8'h6F;
Memory[22675] = 8'h49;
Memory[22674] = 8'h8D;
Memory[22673] = 8'h21;
Memory[22672] = 8'h83;
Memory[22679] = 8'h00;
Memory[22678] = 8'h3B;
Memory[22677] = 8'h2A;
Memory[22676] = 8'h23;
Memory[22683] = 8'h12;
Memory[22682] = 8'h40;
Memory[22681] = 8'h20;
Memory[22680] = 8'h6F;
Memory[22687] = 8'h49;
Memory[22686] = 8'hCD;
Memory[22685] = 8'h21;
Memory[22684] = 8'h83;
Memory[22691] = 8'h00;
Memory[22690] = 8'h3B;
Memory[22689] = 8'h2A;
Memory[22688] = 8'h23;
Memory[22695] = 8'h12;
Memory[22694] = 8'h40;
Memory[22693] = 8'h20;
Memory[22692] = 8'h6F;
Memory[22699] = 8'h4A;
Memory[22698] = 8'h0D;
Memory[22697] = 8'h21;
Memory[22696] = 8'h83;
Memory[22703] = 8'h00;
Memory[22702] = 8'h3B;
Memory[22701] = 8'h2A;
Memory[22700] = 8'h23;
Memory[22707] = 8'h12;
Memory[22706] = 8'h40;
Memory[22705] = 8'h20;
Memory[22704] = 8'h6F;
Memory[22711] = 8'h4A;
Memory[22710] = 8'h4D;
Memory[22709] = 8'h21;
Memory[22708] = 8'h83;
Memory[22715] = 8'h00;
Memory[22714] = 8'h3B;
Memory[22713] = 8'h2A;
Memory[22712] = 8'h23;
Memory[22719] = 8'h12;
Memory[22718] = 8'h40;
Memory[22717] = 8'h20;
Memory[22716] = 8'h6F;
Memory[22723] = 8'h4A;
Memory[22722] = 8'h8D;
Memory[22721] = 8'h21;
Memory[22720] = 8'h83;
Memory[22727] = 8'h00;
Memory[22726] = 8'h3B;
Memory[22725] = 8'h2A;
Memory[22724] = 8'h23;
Memory[22731] = 8'h12;
Memory[22730] = 8'h40;
Memory[22729] = 8'h20;
Memory[22728] = 8'h6F;
Memory[22735] = 8'h4A;
Memory[22734] = 8'hCD;
Memory[22733] = 8'h21;
Memory[22732] = 8'h83;
Memory[22739] = 8'h00;
Memory[22738] = 8'h3B;
Memory[22737] = 8'h2A;
Memory[22736] = 8'h23;
Memory[22743] = 8'h12;
Memory[22742] = 8'h40;
Memory[22741] = 8'h20;
Memory[22740] = 8'h6F;
Memory[22747] = 8'h4B;
Memory[22746] = 8'h0D;
Memory[22745] = 8'h21;
Memory[22744] = 8'h83;
Memory[22751] = 8'h00;
Memory[22750] = 8'h3B;
Memory[22749] = 8'h2A;
Memory[22748] = 8'h23;
Memory[22755] = 8'h12;
Memory[22754] = 8'h40;
Memory[22753] = 8'h20;
Memory[22752] = 8'h6F;
Memory[22759] = 8'h4B;
Memory[22758] = 8'h4D;
Memory[22757] = 8'h21;
Memory[22756] = 8'h83;
Memory[22763] = 8'h00;
Memory[22762] = 8'h3B;
Memory[22761] = 8'h2A;
Memory[22760] = 8'h23;
Memory[22767] = 8'h12;
Memory[22766] = 8'h40;
Memory[22765] = 8'h20;
Memory[22764] = 8'h6F;
Memory[22771] = 8'h4B;
Memory[22770] = 8'h8D;
Memory[22769] = 8'h21;
Memory[22768] = 8'h83;
Memory[22775] = 8'h00;
Memory[22774] = 8'h3B;
Memory[22773] = 8'h2A;
Memory[22772] = 8'h23;
Memory[22779] = 8'h12;
Memory[22778] = 8'h40;
Memory[22777] = 8'h20;
Memory[22776] = 8'h6F;
Memory[22783] = 8'h4B;
Memory[22782] = 8'hCD;
Memory[22781] = 8'h21;
Memory[22780] = 8'h83;
Memory[22787] = 8'h00;
Memory[22786] = 8'h3B;
Memory[22785] = 8'h2A;
Memory[22784] = 8'h23;
Memory[22791] = 8'h12;
Memory[22790] = 8'h40;
Memory[22789] = 8'h20;
Memory[22788] = 8'h6F;
Memory[22795] = 8'h4C;
Memory[22794] = 8'h0D;
Memory[22793] = 8'h21;
Memory[22792] = 8'h83;
Memory[22799] = 8'h00;
Memory[22798] = 8'h3B;
Memory[22797] = 8'h2A;
Memory[22796] = 8'h23;
Memory[22803] = 8'h12;
Memory[22802] = 8'h40;
Memory[22801] = 8'h20;
Memory[22800] = 8'h6F;
Memory[22807] = 8'h4C;
Memory[22806] = 8'h4D;
Memory[22805] = 8'h21;
Memory[22804] = 8'h83;
Memory[22811] = 8'h00;
Memory[22810] = 8'h3B;
Memory[22809] = 8'h2A;
Memory[22808] = 8'h23;
Memory[22815] = 8'h12;
Memory[22814] = 8'h40;
Memory[22813] = 8'h20;
Memory[22812] = 8'h6F;
Memory[22819] = 8'h4C;
Memory[22818] = 8'h8D;
Memory[22817] = 8'h21;
Memory[22816] = 8'h83;
Memory[22823] = 8'h00;
Memory[22822] = 8'h3B;
Memory[22821] = 8'h2A;
Memory[22820] = 8'h23;
Memory[22827] = 8'h12;
Memory[22826] = 8'h40;
Memory[22825] = 8'h20;
Memory[22824] = 8'h6F;
Memory[22831] = 8'h4C;
Memory[22830] = 8'hCD;
Memory[22829] = 8'h21;
Memory[22828] = 8'h83;
Memory[22835] = 8'h00;
Memory[22834] = 8'h3B;
Memory[22833] = 8'h2A;
Memory[22832] = 8'h23;
Memory[22839] = 8'h12;
Memory[22838] = 8'h40;
Memory[22837] = 8'h20;
Memory[22836] = 8'h6F;
Memory[22843] = 8'h4D;
Memory[22842] = 8'h0D;
Memory[22841] = 8'h21;
Memory[22840] = 8'h83;
Memory[22847] = 8'h00;
Memory[22846] = 8'h3B;
Memory[22845] = 8'h2A;
Memory[22844] = 8'h23;
Memory[22851] = 8'h12;
Memory[22850] = 8'h40;
Memory[22849] = 8'h20;
Memory[22848] = 8'h6F;
Memory[22855] = 8'h4D;
Memory[22854] = 8'h4D;
Memory[22853] = 8'h21;
Memory[22852] = 8'h83;
Memory[22859] = 8'h00;
Memory[22858] = 8'h3B;
Memory[22857] = 8'h2A;
Memory[22856] = 8'h23;
Memory[22863] = 8'h12;
Memory[22862] = 8'h40;
Memory[22861] = 8'h20;
Memory[22860] = 8'h6F;
Memory[22867] = 8'h4D;
Memory[22866] = 8'h8D;
Memory[22865] = 8'h21;
Memory[22864] = 8'h83;
Memory[22871] = 8'h00;
Memory[22870] = 8'h3B;
Memory[22869] = 8'h2A;
Memory[22868] = 8'h23;
Memory[22875] = 8'h12;
Memory[22874] = 8'h40;
Memory[22873] = 8'h20;
Memory[22872] = 8'h6F;
Memory[22879] = 8'h4D;
Memory[22878] = 8'hCD;
Memory[22877] = 8'h21;
Memory[22876] = 8'h83;
Memory[22883] = 8'h00;
Memory[22882] = 8'h3B;
Memory[22881] = 8'h2A;
Memory[22880] = 8'h23;
Memory[22887] = 8'h12;
Memory[22886] = 8'h40;
Memory[22885] = 8'h20;
Memory[22884] = 8'h6F;
Memory[22891] = 8'h4E;
Memory[22890] = 8'h0D;
Memory[22889] = 8'h21;
Memory[22888] = 8'h83;
Memory[22895] = 8'h00;
Memory[22894] = 8'h3B;
Memory[22893] = 8'h2A;
Memory[22892] = 8'h23;
Memory[22899] = 8'h12;
Memory[22898] = 8'h40;
Memory[22897] = 8'h20;
Memory[22896] = 8'h6F;
Memory[22903] = 8'h4E;
Memory[22902] = 8'h4D;
Memory[22901] = 8'h21;
Memory[22900] = 8'h83;
Memory[22907] = 8'h00;
Memory[22906] = 8'h3B;
Memory[22905] = 8'h2A;
Memory[22904] = 8'h23;
Memory[22911] = 8'h12;
Memory[22910] = 8'h40;
Memory[22909] = 8'h20;
Memory[22908] = 8'h6F;
Memory[22915] = 8'h4E;
Memory[22914] = 8'h8D;
Memory[22913] = 8'h21;
Memory[22912] = 8'h83;
Memory[22919] = 8'h00;
Memory[22918] = 8'h3B;
Memory[22917] = 8'h2A;
Memory[22916] = 8'h23;
Memory[22923] = 8'h12;
Memory[22922] = 8'h40;
Memory[22921] = 8'h20;
Memory[22920] = 8'h6F;
Memory[22927] = 8'h4E;
Memory[22926] = 8'hCD;
Memory[22925] = 8'h21;
Memory[22924] = 8'h83;
Memory[22931] = 8'h00;
Memory[22930] = 8'h3B;
Memory[22929] = 8'h2A;
Memory[22928] = 8'h23;
Memory[22935] = 8'h12;
Memory[22934] = 8'h40;
Memory[22933] = 8'h20;
Memory[22932] = 8'h6F;
Memory[22939] = 8'h4F;
Memory[22938] = 8'h0D;
Memory[22937] = 8'h21;
Memory[22936] = 8'h83;
Memory[22943] = 8'h00;
Memory[22942] = 8'h3B;
Memory[22941] = 8'h2A;
Memory[22940] = 8'h23;
Memory[22947] = 8'h12;
Memory[22946] = 8'h40;
Memory[22945] = 8'h20;
Memory[22944] = 8'h6F;
Memory[22951] = 8'h4F;
Memory[22950] = 8'h4D;
Memory[22949] = 8'h21;
Memory[22948] = 8'h83;
Memory[22955] = 8'h00;
Memory[22954] = 8'h3B;
Memory[22953] = 8'h2A;
Memory[22952] = 8'h23;
Memory[22959] = 8'h12;
Memory[22958] = 8'h40;
Memory[22957] = 8'h20;
Memory[22956] = 8'h6F;
Memory[22963] = 8'h4F;
Memory[22962] = 8'h8D;
Memory[22961] = 8'h21;
Memory[22960] = 8'h83;
Memory[22967] = 8'h00;
Memory[22966] = 8'h3B;
Memory[22965] = 8'h2A;
Memory[22964] = 8'h23;
Memory[22971] = 8'h12;
Memory[22970] = 8'h40;
Memory[22969] = 8'h20;
Memory[22968] = 8'h6F;
Memory[22975] = 8'h4F;
Memory[22974] = 8'hCD;
Memory[22973] = 8'h21;
Memory[22972] = 8'h83;
Memory[22979] = 8'h00;
Memory[22978] = 8'h3B;
Memory[22977] = 8'h2A;
Memory[22976] = 8'h23;
Memory[22983] = 8'h12;
Memory[22982] = 8'h40;
Memory[22981] = 8'h20;
Memory[22980] = 8'h6F;
Memory[22987] = 8'h50;
Memory[22986] = 8'h0D;
Memory[22985] = 8'h21;
Memory[22984] = 8'h83;
Memory[22991] = 8'h00;
Memory[22990] = 8'h3B;
Memory[22989] = 8'h2A;
Memory[22988] = 8'h23;
Memory[22995] = 8'h12;
Memory[22994] = 8'h40;
Memory[22993] = 8'h20;
Memory[22992] = 8'h6F;
Memory[22999] = 8'h50;
Memory[22998] = 8'h4D;
Memory[22997] = 8'h21;
Memory[22996] = 8'h83;
Memory[23003] = 8'h00;
Memory[23002] = 8'h3B;
Memory[23001] = 8'h2A;
Memory[23000] = 8'h23;
Memory[23007] = 8'h12;
Memory[23006] = 8'h40;
Memory[23005] = 8'h20;
Memory[23004] = 8'h6F;
Memory[23011] = 8'h50;
Memory[23010] = 8'h8D;
Memory[23009] = 8'h21;
Memory[23008] = 8'h83;
Memory[23015] = 8'h00;
Memory[23014] = 8'h3B;
Memory[23013] = 8'h2A;
Memory[23012] = 8'h23;
Memory[23019] = 8'h12;
Memory[23018] = 8'h40;
Memory[23017] = 8'h20;
Memory[23016] = 8'h6F;
Memory[23023] = 8'h50;
Memory[23022] = 8'hCD;
Memory[23021] = 8'h21;
Memory[23020] = 8'h83;
Memory[23027] = 8'h00;
Memory[23026] = 8'h3B;
Memory[23025] = 8'h2A;
Memory[23024] = 8'h23;
Memory[23031] = 8'h12;
Memory[23030] = 8'h40;
Memory[23029] = 8'h20;
Memory[23028] = 8'h6F;
Memory[23035] = 8'h51;
Memory[23034] = 8'h0D;
Memory[23033] = 8'h21;
Memory[23032] = 8'h83;
Memory[23039] = 8'h00;
Memory[23038] = 8'h3B;
Memory[23037] = 8'h2A;
Memory[23036] = 8'h23;
Memory[23043] = 8'h12;
Memory[23042] = 8'h40;
Memory[23041] = 8'h20;
Memory[23040] = 8'h6F;
Memory[23047] = 8'h51;
Memory[23046] = 8'h4D;
Memory[23045] = 8'h21;
Memory[23044] = 8'h83;
Memory[23051] = 8'h00;
Memory[23050] = 8'h3B;
Memory[23049] = 8'h2A;
Memory[23048] = 8'h23;
Memory[23055] = 8'h12;
Memory[23054] = 8'h40;
Memory[23053] = 8'h20;
Memory[23052] = 8'h6F;
Memory[23059] = 8'h51;
Memory[23058] = 8'h8D;
Memory[23057] = 8'h21;
Memory[23056] = 8'h83;
Memory[23063] = 8'h00;
Memory[23062] = 8'h3B;
Memory[23061] = 8'h2A;
Memory[23060] = 8'h23;
Memory[23067] = 8'h12;
Memory[23066] = 8'h40;
Memory[23065] = 8'h20;
Memory[23064] = 8'h6F;
Memory[23071] = 8'h51;
Memory[23070] = 8'hCD;
Memory[23069] = 8'h21;
Memory[23068] = 8'h83;
Memory[23075] = 8'h00;
Memory[23074] = 8'h3B;
Memory[23073] = 8'h2A;
Memory[23072] = 8'h23;
Memory[23079] = 8'h12;
Memory[23078] = 8'h40;
Memory[23077] = 8'h20;
Memory[23076] = 8'h6F;
Memory[23083] = 8'h52;
Memory[23082] = 8'h0D;
Memory[23081] = 8'h21;
Memory[23080] = 8'h83;
Memory[23087] = 8'h00;
Memory[23086] = 8'h3B;
Memory[23085] = 8'h2A;
Memory[23084] = 8'h23;
Memory[23091] = 8'h12;
Memory[23090] = 8'h40;
Memory[23089] = 8'h20;
Memory[23088] = 8'h6F;
Memory[23095] = 8'h52;
Memory[23094] = 8'h4D;
Memory[23093] = 8'h21;
Memory[23092] = 8'h83;
Memory[23099] = 8'h00;
Memory[23098] = 8'h3B;
Memory[23097] = 8'h2A;
Memory[23096] = 8'h23;
Memory[23103] = 8'h12;
Memory[23102] = 8'h40;
Memory[23101] = 8'h20;
Memory[23100] = 8'h6F;
Memory[23107] = 8'h52;
Memory[23106] = 8'h8D;
Memory[23105] = 8'h21;
Memory[23104] = 8'h83;
Memory[23111] = 8'h00;
Memory[23110] = 8'h3B;
Memory[23109] = 8'h2A;
Memory[23108] = 8'h23;
Memory[23115] = 8'h12;
Memory[23114] = 8'h40;
Memory[23113] = 8'h20;
Memory[23112] = 8'h6F;
Memory[23119] = 8'h52;
Memory[23118] = 8'hCD;
Memory[23117] = 8'h21;
Memory[23116] = 8'h83;
Memory[23123] = 8'h00;
Memory[23122] = 8'h3B;
Memory[23121] = 8'h2A;
Memory[23120] = 8'h23;
Memory[23127] = 8'h12;
Memory[23126] = 8'h40;
Memory[23125] = 8'h20;
Memory[23124] = 8'h6F;
Memory[23131] = 8'h53;
Memory[23130] = 8'h0D;
Memory[23129] = 8'h21;
Memory[23128] = 8'h83;
Memory[23135] = 8'h00;
Memory[23134] = 8'h3B;
Memory[23133] = 8'h2A;
Memory[23132] = 8'h23;
Memory[23139] = 8'h12;
Memory[23138] = 8'h40;
Memory[23137] = 8'h20;
Memory[23136] = 8'h6F;
Memory[23143] = 8'h53;
Memory[23142] = 8'h4D;
Memory[23141] = 8'h21;
Memory[23140] = 8'h83;
Memory[23147] = 8'h00;
Memory[23146] = 8'h3B;
Memory[23145] = 8'h2A;
Memory[23144] = 8'h23;
Memory[23151] = 8'h12;
Memory[23150] = 8'h40;
Memory[23149] = 8'h20;
Memory[23148] = 8'h6F;
Memory[23155] = 8'h53;
Memory[23154] = 8'h8D;
Memory[23153] = 8'h21;
Memory[23152] = 8'h83;
Memory[23159] = 8'h00;
Memory[23158] = 8'h3B;
Memory[23157] = 8'h2A;
Memory[23156] = 8'h23;
Memory[23163] = 8'h12;
Memory[23162] = 8'h40;
Memory[23161] = 8'h20;
Memory[23160] = 8'h6F;
Memory[23167] = 8'h53;
Memory[23166] = 8'hCD;
Memory[23165] = 8'h21;
Memory[23164] = 8'h83;
Memory[23171] = 8'h00;
Memory[23170] = 8'h3B;
Memory[23169] = 8'h2A;
Memory[23168] = 8'h23;
Memory[23175] = 8'h12;
Memory[23174] = 8'h40;
Memory[23173] = 8'h20;
Memory[23172] = 8'h6F;
Memory[23179] = 8'h54;
Memory[23178] = 8'h0D;
Memory[23177] = 8'h21;
Memory[23176] = 8'h83;
Memory[23183] = 8'h00;
Memory[23182] = 8'h3B;
Memory[23181] = 8'h2A;
Memory[23180] = 8'h23;
Memory[23187] = 8'h12;
Memory[23186] = 8'h40;
Memory[23185] = 8'h20;
Memory[23184] = 8'h6F;
Memory[23191] = 8'h54;
Memory[23190] = 8'h4D;
Memory[23189] = 8'h21;
Memory[23188] = 8'h83;
Memory[23195] = 8'h00;
Memory[23194] = 8'h3B;
Memory[23193] = 8'h2A;
Memory[23192] = 8'h23;
Memory[23199] = 8'h12;
Memory[23198] = 8'h40;
Memory[23197] = 8'h20;
Memory[23196] = 8'h6F;
Memory[23203] = 8'h54;
Memory[23202] = 8'h8D;
Memory[23201] = 8'h21;
Memory[23200] = 8'h83;
Memory[23207] = 8'h00;
Memory[23206] = 8'h3B;
Memory[23205] = 8'h2A;
Memory[23204] = 8'h23;
Memory[23211] = 8'h12;
Memory[23210] = 8'h40;
Memory[23209] = 8'h20;
Memory[23208] = 8'h6F;
Memory[23215] = 8'h54;
Memory[23214] = 8'hCD;
Memory[23213] = 8'h21;
Memory[23212] = 8'h83;
Memory[23219] = 8'h00;
Memory[23218] = 8'h3B;
Memory[23217] = 8'h2A;
Memory[23216] = 8'h23;
Memory[23223] = 8'h12;
Memory[23222] = 8'h40;
Memory[23221] = 8'h20;
Memory[23220] = 8'h6F;
Memory[23227] = 8'h55;
Memory[23226] = 8'h0D;
Memory[23225] = 8'h21;
Memory[23224] = 8'h83;
Memory[23231] = 8'h00;
Memory[23230] = 8'h3B;
Memory[23229] = 8'h2A;
Memory[23228] = 8'h23;
Memory[23235] = 8'h12;
Memory[23234] = 8'h40;
Memory[23233] = 8'h20;
Memory[23232] = 8'h6F;
Memory[23239] = 8'h55;
Memory[23238] = 8'h4D;
Memory[23237] = 8'h21;
Memory[23236] = 8'h83;
Memory[23243] = 8'h00;
Memory[23242] = 8'h3B;
Memory[23241] = 8'h2A;
Memory[23240] = 8'h23;
Memory[23247] = 8'h12;
Memory[23246] = 8'h40;
Memory[23245] = 8'h20;
Memory[23244] = 8'h6F;
Memory[23251] = 8'h55;
Memory[23250] = 8'h8D;
Memory[23249] = 8'h21;
Memory[23248] = 8'h83;
Memory[23255] = 8'h00;
Memory[23254] = 8'h3B;
Memory[23253] = 8'h2A;
Memory[23252] = 8'h23;
Memory[23259] = 8'h12;
Memory[23258] = 8'h40;
Memory[23257] = 8'h20;
Memory[23256] = 8'h6F;
Memory[23263] = 8'h55;
Memory[23262] = 8'hCD;
Memory[23261] = 8'h21;
Memory[23260] = 8'h83;
Memory[23267] = 8'h00;
Memory[23266] = 8'h3B;
Memory[23265] = 8'h2A;
Memory[23264] = 8'h23;
Memory[23271] = 8'h12;
Memory[23270] = 8'h40;
Memory[23269] = 8'h20;
Memory[23268] = 8'h6F;
Memory[23275] = 8'h56;
Memory[23274] = 8'h0D;
Memory[23273] = 8'h21;
Memory[23272] = 8'h83;
Memory[23279] = 8'h00;
Memory[23278] = 8'h3B;
Memory[23277] = 8'h2A;
Memory[23276] = 8'h23;
Memory[23283] = 8'h12;
Memory[23282] = 8'h40;
Memory[23281] = 8'h20;
Memory[23280] = 8'h6F;
Memory[23287] = 8'h56;
Memory[23286] = 8'h4D;
Memory[23285] = 8'h21;
Memory[23284] = 8'h83;
Memory[23291] = 8'h00;
Memory[23290] = 8'h3B;
Memory[23289] = 8'h2A;
Memory[23288] = 8'h23;
Memory[23295] = 8'h12;
Memory[23294] = 8'h40;
Memory[23293] = 8'h20;
Memory[23292] = 8'h6F;
Memory[23299] = 8'h56;
Memory[23298] = 8'h8D;
Memory[23297] = 8'h21;
Memory[23296] = 8'h83;
Memory[23303] = 8'h00;
Memory[23302] = 8'h3B;
Memory[23301] = 8'h2A;
Memory[23300] = 8'h23;
Memory[23307] = 8'h12;
Memory[23306] = 8'h40;
Memory[23305] = 8'h20;
Memory[23304] = 8'h6F;
Memory[23311] = 8'h56;
Memory[23310] = 8'hCD;
Memory[23309] = 8'h21;
Memory[23308] = 8'h83;
Memory[23315] = 8'h00;
Memory[23314] = 8'h3B;
Memory[23313] = 8'h2A;
Memory[23312] = 8'h23;
Memory[23319] = 8'h12;
Memory[23318] = 8'h40;
Memory[23317] = 8'h20;
Memory[23316] = 8'h6F;
Memory[23323] = 8'h57;
Memory[23322] = 8'h0D;
Memory[23321] = 8'h21;
Memory[23320] = 8'h83;
Memory[23327] = 8'h00;
Memory[23326] = 8'h3B;
Memory[23325] = 8'h2A;
Memory[23324] = 8'h23;
Memory[23331] = 8'h12;
Memory[23330] = 8'h40;
Memory[23329] = 8'h20;
Memory[23328] = 8'h6F;
Memory[23335] = 8'h57;
Memory[23334] = 8'h4D;
Memory[23333] = 8'h21;
Memory[23332] = 8'h83;
Memory[23339] = 8'h00;
Memory[23338] = 8'h3B;
Memory[23337] = 8'h2A;
Memory[23336] = 8'h23;
Memory[23343] = 8'h12;
Memory[23342] = 8'h40;
Memory[23341] = 8'h20;
Memory[23340] = 8'h6F;
Memory[23347] = 8'h57;
Memory[23346] = 8'h8D;
Memory[23345] = 8'h21;
Memory[23344] = 8'h83;
Memory[23351] = 8'h00;
Memory[23350] = 8'h3B;
Memory[23349] = 8'h2A;
Memory[23348] = 8'h23;
Memory[23355] = 8'h12;
Memory[23354] = 8'h40;
Memory[23353] = 8'h20;
Memory[23352] = 8'h6F;
Memory[23359] = 8'h57;
Memory[23358] = 8'hCD;
Memory[23357] = 8'h21;
Memory[23356] = 8'h83;
Memory[23363] = 8'h00;
Memory[23362] = 8'h3B;
Memory[23361] = 8'h2A;
Memory[23360] = 8'h23;
Memory[23367] = 8'h12;
Memory[23366] = 8'h40;
Memory[23365] = 8'h20;
Memory[23364] = 8'h6F;
Memory[23371] = 8'h58;
Memory[23370] = 8'h0D;
Memory[23369] = 8'h21;
Memory[23368] = 8'h83;
Memory[23375] = 8'h00;
Memory[23374] = 8'h3B;
Memory[23373] = 8'h2A;
Memory[23372] = 8'h23;
Memory[23379] = 8'h12;
Memory[23378] = 8'h40;
Memory[23377] = 8'h20;
Memory[23376] = 8'h6F;
Memory[23383] = 8'h58;
Memory[23382] = 8'h4D;
Memory[23381] = 8'h21;
Memory[23380] = 8'h83;
Memory[23387] = 8'h00;
Memory[23386] = 8'h3B;
Memory[23385] = 8'h2A;
Memory[23384] = 8'h23;
Memory[23391] = 8'h12;
Memory[23390] = 8'h40;
Memory[23389] = 8'h20;
Memory[23388] = 8'h6F;
Memory[23395] = 8'h58;
Memory[23394] = 8'h8D;
Memory[23393] = 8'h21;
Memory[23392] = 8'h83;
Memory[23399] = 8'h00;
Memory[23398] = 8'h3B;
Memory[23397] = 8'h2A;
Memory[23396] = 8'h23;
Memory[23403] = 8'h12;
Memory[23402] = 8'h40;
Memory[23401] = 8'h20;
Memory[23400] = 8'h6F;
Memory[23407] = 8'h58;
Memory[23406] = 8'hCD;
Memory[23405] = 8'h21;
Memory[23404] = 8'h83;
Memory[23411] = 8'h00;
Memory[23410] = 8'h3B;
Memory[23409] = 8'h2A;
Memory[23408] = 8'h23;
Memory[23415] = 8'h12;
Memory[23414] = 8'h40;
Memory[23413] = 8'h20;
Memory[23412] = 8'h6F;
Memory[23419] = 8'h59;
Memory[23418] = 8'h0D;
Memory[23417] = 8'h21;
Memory[23416] = 8'h83;
Memory[23423] = 8'h00;
Memory[23422] = 8'h3B;
Memory[23421] = 8'h2A;
Memory[23420] = 8'h23;
Memory[23427] = 8'h12;
Memory[23426] = 8'h40;
Memory[23425] = 8'h20;
Memory[23424] = 8'h6F;
Memory[23431] = 8'h59;
Memory[23430] = 8'h4D;
Memory[23429] = 8'h21;
Memory[23428] = 8'h83;
Memory[23435] = 8'h00;
Memory[23434] = 8'h3B;
Memory[23433] = 8'h2A;
Memory[23432] = 8'h23;
Memory[23439] = 8'h12;
Memory[23438] = 8'h40;
Memory[23437] = 8'h20;
Memory[23436] = 8'h6F;
Memory[23443] = 8'h59;
Memory[23442] = 8'h8D;
Memory[23441] = 8'h21;
Memory[23440] = 8'h83;
Memory[23447] = 8'h00;
Memory[23446] = 8'h3B;
Memory[23445] = 8'h2A;
Memory[23444] = 8'h23;
Memory[23451] = 8'h12;
Memory[23450] = 8'h40;
Memory[23449] = 8'h20;
Memory[23448] = 8'h6F;
Memory[23455] = 8'h59;
Memory[23454] = 8'hCD;
Memory[23453] = 8'h21;
Memory[23452] = 8'h83;
Memory[23459] = 8'h00;
Memory[23458] = 8'h3B;
Memory[23457] = 8'h2A;
Memory[23456] = 8'h23;
Memory[23463] = 8'h12;
Memory[23462] = 8'h40;
Memory[23461] = 8'h20;
Memory[23460] = 8'h6F;
Memory[23467] = 8'h5A;
Memory[23466] = 8'h0D;
Memory[23465] = 8'h21;
Memory[23464] = 8'h83;
Memory[23471] = 8'h00;
Memory[23470] = 8'h3B;
Memory[23469] = 8'h2A;
Memory[23468] = 8'h23;
Memory[23475] = 8'h12;
Memory[23474] = 8'h40;
Memory[23473] = 8'h20;
Memory[23472] = 8'h6F;
Memory[23479] = 8'h5A;
Memory[23478] = 8'h4D;
Memory[23477] = 8'h21;
Memory[23476] = 8'h83;
Memory[23483] = 8'h00;
Memory[23482] = 8'h3B;
Memory[23481] = 8'h2A;
Memory[23480] = 8'h23;
Memory[23487] = 8'h12;
Memory[23486] = 8'h40;
Memory[23485] = 8'h20;
Memory[23484] = 8'h6F;
Memory[23491] = 8'h5A;
Memory[23490] = 8'h8D;
Memory[23489] = 8'h21;
Memory[23488] = 8'h83;
Memory[23495] = 8'h00;
Memory[23494] = 8'h3B;
Memory[23493] = 8'h2A;
Memory[23492] = 8'h23;
Memory[23499] = 8'h12;
Memory[23498] = 8'h40;
Memory[23497] = 8'h20;
Memory[23496] = 8'h6F;
Memory[23503] = 8'h5A;
Memory[23502] = 8'hCD;
Memory[23501] = 8'h21;
Memory[23500] = 8'h83;
Memory[23507] = 8'h00;
Memory[23506] = 8'h3B;
Memory[23505] = 8'h2A;
Memory[23504] = 8'h23;
Memory[23511] = 8'h12;
Memory[23510] = 8'h40;
Memory[23509] = 8'h20;
Memory[23508] = 8'h6F;
Memory[23515] = 8'h5B;
Memory[23514] = 8'h0D;
Memory[23513] = 8'h21;
Memory[23512] = 8'h83;
Memory[23519] = 8'h00;
Memory[23518] = 8'h3B;
Memory[23517] = 8'h2A;
Memory[23516] = 8'h23;
Memory[23523] = 8'h12;
Memory[23522] = 8'h40;
Memory[23521] = 8'h20;
Memory[23520] = 8'h6F;
Memory[23527] = 8'h5B;
Memory[23526] = 8'h4D;
Memory[23525] = 8'h21;
Memory[23524] = 8'h83;
Memory[23531] = 8'h00;
Memory[23530] = 8'h3B;
Memory[23529] = 8'h2A;
Memory[23528] = 8'h23;
Memory[23535] = 8'h12;
Memory[23534] = 8'h40;
Memory[23533] = 8'h20;
Memory[23532] = 8'h6F;
Memory[23539] = 8'h5B;
Memory[23538] = 8'h8D;
Memory[23537] = 8'h21;
Memory[23536] = 8'h83;
Memory[23543] = 8'h00;
Memory[23542] = 8'h3B;
Memory[23541] = 8'h2A;
Memory[23540] = 8'h23;
Memory[23547] = 8'h12;
Memory[23546] = 8'h40;
Memory[23545] = 8'h20;
Memory[23544] = 8'h6F;
Memory[23551] = 8'h5B;
Memory[23550] = 8'hCD;
Memory[23549] = 8'h21;
Memory[23548] = 8'h83;
Memory[23555] = 8'h00;
Memory[23554] = 8'h3B;
Memory[23553] = 8'h2A;
Memory[23552] = 8'h23;
Memory[23559] = 8'h12;
Memory[23558] = 8'h40;
Memory[23557] = 8'h20;
Memory[23556] = 8'h6F;
Memory[23563] = 8'h5C;
Memory[23562] = 8'h0D;
Memory[23561] = 8'h21;
Memory[23560] = 8'h83;
Memory[23567] = 8'h00;
Memory[23566] = 8'h3B;
Memory[23565] = 8'h2A;
Memory[23564] = 8'h23;
Memory[23571] = 8'h12;
Memory[23570] = 8'h40;
Memory[23569] = 8'h20;
Memory[23568] = 8'h6F;
Memory[23575] = 8'h5C;
Memory[23574] = 8'h4D;
Memory[23573] = 8'h21;
Memory[23572] = 8'h83;
Memory[23579] = 8'h00;
Memory[23578] = 8'h3B;
Memory[23577] = 8'h2A;
Memory[23576] = 8'h23;
Memory[23583] = 8'h12;
Memory[23582] = 8'h40;
Memory[23581] = 8'h20;
Memory[23580] = 8'h6F;
Memory[23587] = 8'h5C;
Memory[23586] = 8'h8D;
Memory[23585] = 8'h21;
Memory[23584] = 8'h83;
Memory[23591] = 8'h00;
Memory[23590] = 8'h3B;
Memory[23589] = 8'h2A;
Memory[23588] = 8'h23;
Memory[23595] = 8'h12;
Memory[23594] = 8'h40;
Memory[23593] = 8'h20;
Memory[23592] = 8'h6F;
Memory[23599] = 8'h5C;
Memory[23598] = 8'hCD;
Memory[23597] = 8'h21;
Memory[23596] = 8'h83;
Memory[23603] = 8'h00;
Memory[23602] = 8'h3B;
Memory[23601] = 8'h2A;
Memory[23600] = 8'h23;
Memory[23607] = 8'h12;
Memory[23606] = 8'h40;
Memory[23605] = 8'h20;
Memory[23604] = 8'h6F;
Memory[23611] = 8'h5D;
Memory[23610] = 8'h0D;
Memory[23609] = 8'h21;
Memory[23608] = 8'h83;
Memory[23615] = 8'h00;
Memory[23614] = 8'h3B;
Memory[23613] = 8'h2A;
Memory[23612] = 8'h23;
Memory[23619] = 8'h12;
Memory[23618] = 8'h40;
Memory[23617] = 8'h20;
Memory[23616] = 8'h6F;
Memory[23623] = 8'h5D;
Memory[23622] = 8'h4D;
Memory[23621] = 8'h21;
Memory[23620] = 8'h83;
Memory[23627] = 8'h00;
Memory[23626] = 8'h3B;
Memory[23625] = 8'h2A;
Memory[23624] = 8'h23;
Memory[23631] = 8'h12;
Memory[23630] = 8'h40;
Memory[23629] = 8'h20;
Memory[23628] = 8'h6F;
Memory[23635] = 8'h5D;
Memory[23634] = 8'h8D;
Memory[23633] = 8'h21;
Memory[23632] = 8'h83;
Memory[23639] = 8'h00;
Memory[23638] = 8'h3B;
Memory[23637] = 8'h2A;
Memory[23636] = 8'h23;
Memory[23643] = 8'h12;
Memory[23642] = 8'h40;
Memory[23641] = 8'h20;
Memory[23640] = 8'h6F;
Memory[23647] = 8'h5D;
Memory[23646] = 8'hCD;
Memory[23645] = 8'h21;
Memory[23644] = 8'h83;
Memory[23651] = 8'h00;
Memory[23650] = 8'h3B;
Memory[23649] = 8'h2A;
Memory[23648] = 8'h23;
Memory[23655] = 8'h12;
Memory[23654] = 8'h40;
Memory[23653] = 8'h20;
Memory[23652] = 8'h6F;
Memory[23659] = 8'h5E;
Memory[23658] = 8'h0D;
Memory[23657] = 8'h21;
Memory[23656] = 8'h83;
Memory[23663] = 8'h00;
Memory[23662] = 8'h3B;
Memory[23661] = 8'h2A;
Memory[23660] = 8'h23;
Memory[23667] = 8'h12;
Memory[23666] = 8'h40;
Memory[23665] = 8'h20;
Memory[23664] = 8'h6F;
Memory[23671] = 8'h5E;
Memory[23670] = 8'h4D;
Memory[23669] = 8'h21;
Memory[23668] = 8'h83;
Memory[23675] = 8'h00;
Memory[23674] = 8'h3B;
Memory[23673] = 8'h2A;
Memory[23672] = 8'h23;
Memory[23679] = 8'h12;
Memory[23678] = 8'h40;
Memory[23677] = 8'h20;
Memory[23676] = 8'h6F;
Memory[23683] = 8'h5E;
Memory[23682] = 8'h8D;
Memory[23681] = 8'h21;
Memory[23680] = 8'h83;
Memory[23687] = 8'h00;
Memory[23686] = 8'h3B;
Memory[23685] = 8'h2A;
Memory[23684] = 8'h23;
Memory[23691] = 8'h12;
Memory[23690] = 8'h40;
Memory[23689] = 8'h20;
Memory[23688] = 8'h6F;
Memory[23695] = 8'h5E;
Memory[23694] = 8'hCD;
Memory[23693] = 8'h21;
Memory[23692] = 8'h83;
Memory[23699] = 8'h00;
Memory[23698] = 8'h3B;
Memory[23697] = 8'h2A;
Memory[23696] = 8'h23;
Memory[23703] = 8'h12;
Memory[23702] = 8'h40;
Memory[23701] = 8'h20;
Memory[23700] = 8'h6F;
Memory[23707] = 8'h5F;
Memory[23706] = 8'h0D;
Memory[23705] = 8'h21;
Memory[23704] = 8'h83;
Memory[23711] = 8'h00;
Memory[23710] = 8'h3B;
Memory[23709] = 8'h2A;
Memory[23708] = 8'h23;
Memory[23715] = 8'h12;
Memory[23714] = 8'h40;
Memory[23713] = 8'h20;
Memory[23712] = 8'h6F;
Memory[23719] = 8'h5F;
Memory[23718] = 8'h4D;
Memory[23717] = 8'h21;
Memory[23716] = 8'h83;
Memory[23723] = 8'h00;
Memory[23722] = 8'h3B;
Memory[23721] = 8'h2A;
Memory[23720] = 8'h23;
Memory[23727] = 8'h12;
Memory[23726] = 8'h40;
Memory[23725] = 8'h20;
Memory[23724] = 8'h6F;
Memory[23731] = 8'h5F;
Memory[23730] = 8'h8D;
Memory[23729] = 8'h21;
Memory[23728] = 8'h83;
Memory[23735] = 8'h00;
Memory[23734] = 8'h3B;
Memory[23733] = 8'h2A;
Memory[23732] = 8'h23;
Memory[23739] = 8'h12;
Memory[23738] = 8'h40;
Memory[23737] = 8'h20;
Memory[23736] = 8'h6F;
Memory[23743] = 8'h5F;
Memory[23742] = 8'hCD;
Memory[23741] = 8'h21;
Memory[23740] = 8'h83;
Memory[23747] = 8'h00;
Memory[23746] = 8'h3B;
Memory[23745] = 8'h2A;
Memory[23744] = 8'h23;
Memory[23751] = 8'h12;
Memory[23750] = 8'h40;
Memory[23749] = 8'h20;
Memory[23748] = 8'h6F;
Memory[23755] = 8'h60;
Memory[23754] = 8'h0D;
Memory[23753] = 8'h21;
Memory[23752] = 8'h83;
Memory[23759] = 8'h00;
Memory[23758] = 8'h3B;
Memory[23757] = 8'h2A;
Memory[23756] = 8'h23;
Memory[23763] = 8'h12;
Memory[23762] = 8'h40;
Memory[23761] = 8'h20;
Memory[23760] = 8'h6F;
Memory[23767] = 8'h60;
Memory[23766] = 8'h4D;
Memory[23765] = 8'h21;
Memory[23764] = 8'h83;
Memory[23771] = 8'h00;
Memory[23770] = 8'h3B;
Memory[23769] = 8'h2A;
Memory[23768] = 8'h23;
Memory[23775] = 8'h12;
Memory[23774] = 8'h40;
Memory[23773] = 8'h20;
Memory[23772] = 8'h6F;
Memory[23779] = 8'h60;
Memory[23778] = 8'h8D;
Memory[23777] = 8'h21;
Memory[23776] = 8'h83;
Memory[23783] = 8'h00;
Memory[23782] = 8'h3B;
Memory[23781] = 8'h2A;
Memory[23780] = 8'h23;
Memory[23787] = 8'h12;
Memory[23786] = 8'h40;
Memory[23785] = 8'h20;
Memory[23784] = 8'h6F;
Memory[23791] = 8'h60;
Memory[23790] = 8'hCD;
Memory[23789] = 8'h21;
Memory[23788] = 8'h83;
Memory[23795] = 8'h00;
Memory[23794] = 8'h3B;
Memory[23793] = 8'h2A;
Memory[23792] = 8'h23;
Memory[23799] = 8'h12;
Memory[23798] = 8'h40;
Memory[23797] = 8'h20;
Memory[23796] = 8'h6F;
Memory[23803] = 8'h61;
Memory[23802] = 8'h0D;
Memory[23801] = 8'h21;
Memory[23800] = 8'h83;
Memory[23807] = 8'h00;
Memory[23806] = 8'h3B;
Memory[23805] = 8'h2A;
Memory[23804] = 8'h23;
Memory[23811] = 8'h12;
Memory[23810] = 8'h40;
Memory[23809] = 8'h20;
Memory[23808] = 8'h6F;
Memory[23815] = 8'h61;
Memory[23814] = 8'h4D;
Memory[23813] = 8'h21;
Memory[23812] = 8'h83;
Memory[23819] = 8'h00;
Memory[23818] = 8'h3B;
Memory[23817] = 8'h2A;
Memory[23816] = 8'h23;
Memory[23823] = 8'h12;
Memory[23822] = 8'h40;
Memory[23821] = 8'h20;
Memory[23820] = 8'h6F;
Memory[23827] = 8'h61;
Memory[23826] = 8'h8D;
Memory[23825] = 8'h21;
Memory[23824] = 8'h83;
Memory[23831] = 8'h00;
Memory[23830] = 8'h3B;
Memory[23829] = 8'h2A;
Memory[23828] = 8'h23;
Memory[23835] = 8'h12;
Memory[23834] = 8'h40;
Memory[23833] = 8'h20;
Memory[23832] = 8'h6F;
Memory[23839] = 8'h61;
Memory[23838] = 8'hCD;
Memory[23837] = 8'h21;
Memory[23836] = 8'h83;
Memory[23843] = 8'h00;
Memory[23842] = 8'h3B;
Memory[23841] = 8'h2A;
Memory[23840] = 8'h23;
Memory[23847] = 8'h12;
Memory[23846] = 8'h40;
Memory[23845] = 8'h20;
Memory[23844] = 8'h6F;
Memory[23851] = 8'h62;
Memory[23850] = 8'h0D;
Memory[23849] = 8'h21;
Memory[23848] = 8'h83;
Memory[23855] = 8'h00;
Memory[23854] = 8'h3B;
Memory[23853] = 8'h2A;
Memory[23852] = 8'h23;
Memory[23859] = 8'h12;
Memory[23858] = 8'h40;
Memory[23857] = 8'h20;
Memory[23856] = 8'h6F;
Memory[23863] = 8'h62;
Memory[23862] = 8'h4D;
Memory[23861] = 8'h21;
Memory[23860] = 8'h83;
Memory[23867] = 8'h00;
Memory[23866] = 8'h3B;
Memory[23865] = 8'h2A;
Memory[23864] = 8'h23;
Memory[23871] = 8'h12;
Memory[23870] = 8'h40;
Memory[23869] = 8'h20;
Memory[23868] = 8'h6F;
Memory[23875] = 8'h62;
Memory[23874] = 8'h8D;
Memory[23873] = 8'h21;
Memory[23872] = 8'h83;
Memory[23879] = 8'h00;
Memory[23878] = 8'h3B;
Memory[23877] = 8'h2A;
Memory[23876] = 8'h23;
Memory[23883] = 8'h12;
Memory[23882] = 8'h40;
Memory[23881] = 8'h20;
Memory[23880] = 8'h6F;
Memory[23887] = 8'h62;
Memory[23886] = 8'hCD;
Memory[23885] = 8'h21;
Memory[23884] = 8'h83;
Memory[23891] = 8'h00;
Memory[23890] = 8'h3B;
Memory[23889] = 8'h2A;
Memory[23888] = 8'h23;
Memory[23895] = 8'h12;
Memory[23894] = 8'h40;
Memory[23893] = 8'h20;
Memory[23892] = 8'h6F;
Memory[23899] = 8'h63;
Memory[23898] = 8'h0D;
Memory[23897] = 8'h21;
Memory[23896] = 8'h83;
Memory[23903] = 8'h00;
Memory[23902] = 8'h3B;
Memory[23901] = 8'h2A;
Memory[23900] = 8'h23;
Memory[23907] = 8'h12;
Memory[23906] = 8'h40;
Memory[23905] = 8'h20;
Memory[23904] = 8'h6F;
Memory[23911] = 8'h63;
Memory[23910] = 8'h4D;
Memory[23909] = 8'h21;
Memory[23908] = 8'h83;
Memory[23915] = 8'h00;
Memory[23914] = 8'h3B;
Memory[23913] = 8'h2A;
Memory[23912] = 8'h23;
Memory[23919] = 8'h12;
Memory[23918] = 8'h40;
Memory[23917] = 8'h20;
Memory[23916] = 8'h6F;
Memory[23923] = 8'h63;
Memory[23922] = 8'h8D;
Memory[23921] = 8'h21;
Memory[23920] = 8'h83;
Memory[23927] = 8'h00;
Memory[23926] = 8'h3B;
Memory[23925] = 8'h2A;
Memory[23924] = 8'h23;
Memory[23931] = 8'h12;
Memory[23930] = 8'h40;
Memory[23929] = 8'h20;
Memory[23928] = 8'h6F;
Memory[23935] = 8'h63;
Memory[23934] = 8'hCD;
Memory[23933] = 8'h21;
Memory[23932] = 8'h83;
Memory[23939] = 8'h00;
Memory[23938] = 8'h3B;
Memory[23937] = 8'h2A;
Memory[23936] = 8'h23;
Memory[23943] = 8'h12;
Memory[23942] = 8'h40;
Memory[23941] = 8'h20;
Memory[23940] = 8'h6F;
Memory[23947] = 8'h64;
Memory[23946] = 8'h0D;
Memory[23945] = 8'h21;
Memory[23944] = 8'h83;
Memory[23951] = 8'h00;
Memory[23950] = 8'h3B;
Memory[23949] = 8'h2A;
Memory[23948] = 8'h23;
Memory[23955] = 8'h12;
Memory[23954] = 8'h40;
Memory[23953] = 8'h20;
Memory[23952] = 8'h6F;
Memory[23959] = 8'h64;
Memory[23958] = 8'h4D;
Memory[23957] = 8'h21;
Memory[23956] = 8'h83;
Memory[23963] = 8'h00;
Memory[23962] = 8'h3B;
Memory[23961] = 8'h2A;
Memory[23960] = 8'h23;
Memory[23967] = 8'h12;
Memory[23966] = 8'h40;
Memory[23965] = 8'h20;
Memory[23964] = 8'h6F;
Memory[23971] = 8'h64;
Memory[23970] = 8'h8D;
Memory[23969] = 8'h21;
Memory[23968] = 8'h83;
Memory[23975] = 8'h00;
Memory[23974] = 8'h3B;
Memory[23973] = 8'h2A;
Memory[23972] = 8'h23;
Memory[23979] = 8'h12;
Memory[23978] = 8'h40;
Memory[23977] = 8'h20;
Memory[23976] = 8'h6F;
Memory[23983] = 8'h64;
Memory[23982] = 8'hCD;
Memory[23981] = 8'h21;
Memory[23980] = 8'h83;
Memory[23987] = 8'h00;
Memory[23986] = 8'h3B;
Memory[23985] = 8'h2A;
Memory[23984] = 8'h23;
Memory[23991] = 8'h12;
Memory[23990] = 8'h40;
Memory[23989] = 8'h20;
Memory[23988] = 8'h6F;
Memory[23995] = 8'h65;
Memory[23994] = 8'h0D;
Memory[23993] = 8'h21;
Memory[23992] = 8'h83;
Memory[23999] = 8'h00;
Memory[23998] = 8'h3B;
Memory[23997] = 8'h2A;
Memory[23996] = 8'h23;
Memory[24003] = 8'h12;
Memory[24002] = 8'h40;
Memory[24001] = 8'h20;
Memory[24000] = 8'h6F;
Memory[24007] = 8'h65;
Memory[24006] = 8'h4D;
Memory[24005] = 8'h21;
Memory[24004] = 8'h83;
Memory[24011] = 8'h00;
Memory[24010] = 8'h3B;
Memory[24009] = 8'h2A;
Memory[24008] = 8'h23;
Memory[24015] = 8'h12;
Memory[24014] = 8'h40;
Memory[24013] = 8'h20;
Memory[24012] = 8'h6F;
Memory[24019] = 8'h65;
Memory[24018] = 8'h8D;
Memory[24017] = 8'h21;
Memory[24016] = 8'h83;
Memory[24023] = 8'h00;
Memory[24022] = 8'h3B;
Memory[24021] = 8'h2A;
Memory[24020] = 8'h23;
Memory[24027] = 8'h12;
Memory[24026] = 8'h40;
Memory[24025] = 8'h20;
Memory[24024] = 8'h6F;
Memory[24031] = 8'h65;
Memory[24030] = 8'hCD;
Memory[24029] = 8'h21;
Memory[24028] = 8'h83;
Memory[24035] = 8'h00;
Memory[24034] = 8'h3B;
Memory[24033] = 8'h2A;
Memory[24032] = 8'h23;
Memory[24039] = 8'h12;
Memory[24038] = 8'h40;
Memory[24037] = 8'h20;
Memory[24036] = 8'h6F;
Memory[24043] = 8'h66;
Memory[24042] = 8'h0D;
Memory[24041] = 8'h21;
Memory[24040] = 8'h83;
Memory[24047] = 8'h00;
Memory[24046] = 8'h3B;
Memory[24045] = 8'h2A;
Memory[24044] = 8'h23;
Memory[24051] = 8'h12;
Memory[24050] = 8'h40;
Memory[24049] = 8'h20;
Memory[24048] = 8'h6F;
Memory[24055] = 8'h66;
Memory[24054] = 8'h4D;
Memory[24053] = 8'h21;
Memory[24052] = 8'h83;
Memory[24059] = 8'h00;
Memory[24058] = 8'h3B;
Memory[24057] = 8'h2A;
Memory[24056] = 8'h23;
Memory[24063] = 8'h12;
Memory[24062] = 8'h40;
Memory[24061] = 8'h20;
Memory[24060] = 8'h6F;
Memory[24067] = 8'h66;
Memory[24066] = 8'h8D;
Memory[24065] = 8'h21;
Memory[24064] = 8'h83;
Memory[24071] = 8'h00;
Memory[24070] = 8'h3B;
Memory[24069] = 8'h2A;
Memory[24068] = 8'h23;
Memory[24075] = 8'h12;
Memory[24074] = 8'h40;
Memory[24073] = 8'h20;
Memory[24072] = 8'h6F;
Memory[24079] = 8'h66;
Memory[24078] = 8'hCD;
Memory[24077] = 8'h21;
Memory[24076] = 8'h83;
Memory[24083] = 8'h00;
Memory[24082] = 8'h3B;
Memory[24081] = 8'h2A;
Memory[24080] = 8'h23;
Memory[24087] = 8'h12;
Memory[24086] = 8'h40;
Memory[24085] = 8'h20;
Memory[24084] = 8'h6F;
Memory[24091] = 8'h67;
Memory[24090] = 8'h0D;
Memory[24089] = 8'h21;
Memory[24088] = 8'h83;
Memory[24095] = 8'h00;
Memory[24094] = 8'h3B;
Memory[24093] = 8'h2A;
Memory[24092] = 8'h23;
Memory[24099] = 8'h12;
Memory[24098] = 8'h40;
Memory[24097] = 8'h20;
Memory[24096] = 8'h6F;
Memory[24103] = 8'h67;
Memory[24102] = 8'h4D;
Memory[24101] = 8'h21;
Memory[24100] = 8'h83;
Memory[24107] = 8'h00;
Memory[24106] = 8'h3B;
Memory[24105] = 8'h2A;
Memory[24104] = 8'h23;
Memory[24111] = 8'h12;
Memory[24110] = 8'h40;
Memory[24109] = 8'h20;
Memory[24108] = 8'h6F;
Memory[24115] = 8'h67;
Memory[24114] = 8'h8D;
Memory[24113] = 8'h21;
Memory[24112] = 8'h83;
Memory[24119] = 8'h00;
Memory[24118] = 8'h3B;
Memory[24117] = 8'h2A;
Memory[24116] = 8'h23;
Memory[24123] = 8'h12;
Memory[24122] = 8'h40;
Memory[24121] = 8'h20;
Memory[24120] = 8'h6F;
Memory[24127] = 8'h67;
Memory[24126] = 8'hCD;
Memory[24125] = 8'h21;
Memory[24124] = 8'h83;
Memory[24131] = 8'h00;
Memory[24130] = 8'h3B;
Memory[24129] = 8'h2A;
Memory[24128] = 8'h23;
Memory[24135] = 8'h12;
Memory[24134] = 8'h40;
Memory[24133] = 8'h20;
Memory[24132] = 8'h6F;
Memory[24139] = 8'h68;
Memory[24138] = 8'h0D;
Memory[24137] = 8'h21;
Memory[24136] = 8'h83;
Memory[24143] = 8'h00;
Memory[24142] = 8'h3B;
Memory[24141] = 8'h2A;
Memory[24140] = 8'h23;
Memory[24147] = 8'h12;
Memory[24146] = 8'h40;
Memory[24145] = 8'h20;
Memory[24144] = 8'h6F;
Memory[24151] = 8'h68;
Memory[24150] = 8'h4D;
Memory[24149] = 8'h21;
Memory[24148] = 8'h83;
Memory[24155] = 8'h00;
Memory[24154] = 8'h3B;
Memory[24153] = 8'h2A;
Memory[24152] = 8'h23;
Memory[24159] = 8'h12;
Memory[24158] = 8'h40;
Memory[24157] = 8'h20;
Memory[24156] = 8'h6F;
Memory[24163] = 8'h68;
Memory[24162] = 8'h8D;
Memory[24161] = 8'h21;
Memory[24160] = 8'h83;
Memory[24167] = 8'h00;
Memory[24166] = 8'h3B;
Memory[24165] = 8'h2A;
Memory[24164] = 8'h23;
Memory[24171] = 8'h12;
Memory[24170] = 8'h40;
Memory[24169] = 8'h20;
Memory[24168] = 8'h6F;
Memory[24175] = 8'h68;
Memory[24174] = 8'hCD;
Memory[24173] = 8'h21;
Memory[24172] = 8'h83;
Memory[24179] = 8'h00;
Memory[24178] = 8'h3B;
Memory[24177] = 8'h2A;
Memory[24176] = 8'h23;
Memory[24183] = 8'h12;
Memory[24182] = 8'h40;
Memory[24181] = 8'h20;
Memory[24180] = 8'h6F;
Memory[24187] = 8'h69;
Memory[24186] = 8'h0D;
Memory[24185] = 8'h21;
Memory[24184] = 8'h83;
Memory[24191] = 8'h00;
Memory[24190] = 8'h3B;
Memory[24189] = 8'h2A;
Memory[24188] = 8'h23;
Memory[24195] = 8'h12;
Memory[24194] = 8'h40;
Memory[24193] = 8'h20;
Memory[24192] = 8'h6F;
Memory[24199] = 8'h69;
Memory[24198] = 8'h4D;
Memory[24197] = 8'h21;
Memory[24196] = 8'h83;
Memory[24203] = 8'h00;
Memory[24202] = 8'h3B;
Memory[24201] = 8'h2A;
Memory[24200] = 8'h23;
Memory[24207] = 8'h12;
Memory[24206] = 8'h40;
Memory[24205] = 8'h20;
Memory[24204] = 8'h6F;
Memory[24211] = 8'h69;
Memory[24210] = 8'h8D;
Memory[24209] = 8'h21;
Memory[24208] = 8'h83;
Memory[24215] = 8'h00;
Memory[24214] = 8'h3B;
Memory[24213] = 8'h2A;
Memory[24212] = 8'h23;
Memory[24219] = 8'h12;
Memory[24218] = 8'h40;
Memory[24217] = 8'h20;
Memory[24216] = 8'h6F;
Memory[24223] = 8'h69;
Memory[24222] = 8'hCD;
Memory[24221] = 8'h21;
Memory[24220] = 8'h83;
Memory[24227] = 8'h00;
Memory[24226] = 8'h3B;
Memory[24225] = 8'h2A;
Memory[24224] = 8'h23;
Memory[24231] = 8'h12;
Memory[24230] = 8'h40;
Memory[24229] = 8'h20;
Memory[24228] = 8'h6F;
Memory[24235] = 8'h6A;
Memory[24234] = 8'h0D;
Memory[24233] = 8'h21;
Memory[24232] = 8'h83;
Memory[24239] = 8'h00;
Memory[24238] = 8'h3B;
Memory[24237] = 8'h2A;
Memory[24236] = 8'h23;
Memory[24243] = 8'h12;
Memory[24242] = 8'h40;
Memory[24241] = 8'h20;
Memory[24240] = 8'h6F;
Memory[24247] = 8'h6A;
Memory[24246] = 8'h4D;
Memory[24245] = 8'h21;
Memory[24244] = 8'h83;
Memory[24251] = 8'h00;
Memory[24250] = 8'h3B;
Memory[24249] = 8'h2A;
Memory[24248] = 8'h23;
Memory[24255] = 8'h12;
Memory[24254] = 8'h40;
Memory[24253] = 8'h20;
Memory[24252] = 8'h6F;
Memory[24259] = 8'h6A;
Memory[24258] = 8'h8D;
Memory[24257] = 8'h21;
Memory[24256] = 8'h83;
Memory[24263] = 8'h00;
Memory[24262] = 8'h3B;
Memory[24261] = 8'h2A;
Memory[24260] = 8'h23;
Memory[24267] = 8'h12;
Memory[24266] = 8'h40;
Memory[24265] = 8'h20;
Memory[24264] = 8'h6F;
Memory[24271] = 8'h6A;
Memory[24270] = 8'hCD;
Memory[24269] = 8'h21;
Memory[24268] = 8'h83;
Memory[24275] = 8'h00;
Memory[24274] = 8'h3B;
Memory[24273] = 8'h2A;
Memory[24272] = 8'h23;
Memory[24279] = 8'h12;
Memory[24278] = 8'h40;
Memory[24277] = 8'h20;
Memory[24276] = 8'h6F;
Memory[24283] = 8'h6B;
Memory[24282] = 8'h0D;
Memory[24281] = 8'h21;
Memory[24280] = 8'h83;
Memory[24287] = 8'h00;
Memory[24286] = 8'h3B;
Memory[24285] = 8'h2A;
Memory[24284] = 8'h23;
Memory[24291] = 8'h12;
Memory[24290] = 8'h40;
Memory[24289] = 8'h20;
Memory[24288] = 8'h6F;
Memory[24295] = 8'h6B;
Memory[24294] = 8'h4D;
Memory[24293] = 8'h21;
Memory[24292] = 8'h83;
Memory[24299] = 8'h00;
Memory[24298] = 8'h3B;
Memory[24297] = 8'h2A;
Memory[24296] = 8'h23;
Memory[24303] = 8'h12;
Memory[24302] = 8'h40;
Memory[24301] = 8'h20;
Memory[24300] = 8'h6F;
Memory[24307] = 8'h6B;
Memory[24306] = 8'h8D;
Memory[24305] = 8'h21;
Memory[24304] = 8'h83;
Memory[24311] = 8'h00;
Memory[24310] = 8'h3B;
Memory[24309] = 8'h2A;
Memory[24308] = 8'h23;
Memory[24315] = 8'h12;
Memory[24314] = 8'h40;
Memory[24313] = 8'h20;
Memory[24312] = 8'h6F;
Memory[24319] = 8'h6B;
Memory[24318] = 8'hCD;
Memory[24317] = 8'h21;
Memory[24316] = 8'h83;
Memory[24323] = 8'h00;
Memory[24322] = 8'h3B;
Memory[24321] = 8'h2A;
Memory[24320] = 8'h23;
Memory[24327] = 8'h12;
Memory[24326] = 8'h40;
Memory[24325] = 8'h20;
Memory[24324] = 8'h6F;
Memory[24331] = 8'h6C;
Memory[24330] = 8'h0D;
Memory[24329] = 8'h21;
Memory[24328] = 8'h83;
Memory[24335] = 8'h00;
Memory[24334] = 8'h3B;
Memory[24333] = 8'h2A;
Memory[24332] = 8'h23;
Memory[24339] = 8'h12;
Memory[24338] = 8'h40;
Memory[24337] = 8'h20;
Memory[24336] = 8'h6F;
Memory[24343] = 8'h6C;
Memory[24342] = 8'h4D;
Memory[24341] = 8'h21;
Memory[24340] = 8'h83;
Memory[24347] = 8'h00;
Memory[24346] = 8'h3B;
Memory[24345] = 8'h2A;
Memory[24344] = 8'h23;
Memory[24351] = 8'h12;
Memory[24350] = 8'h40;
Memory[24349] = 8'h20;
Memory[24348] = 8'h6F;
Memory[24355] = 8'h6C;
Memory[24354] = 8'h8D;
Memory[24353] = 8'h21;
Memory[24352] = 8'h83;
Memory[24359] = 8'h00;
Memory[24358] = 8'h3B;
Memory[24357] = 8'h2A;
Memory[24356] = 8'h23;
Memory[24363] = 8'h12;
Memory[24362] = 8'h40;
Memory[24361] = 8'h20;
Memory[24360] = 8'h6F;
Memory[24367] = 8'h6C;
Memory[24366] = 8'hCD;
Memory[24365] = 8'h21;
Memory[24364] = 8'h83;
Memory[24371] = 8'h00;
Memory[24370] = 8'h3B;
Memory[24369] = 8'h2A;
Memory[24368] = 8'h23;
Memory[24375] = 8'h12;
Memory[24374] = 8'h40;
Memory[24373] = 8'h20;
Memory[24372] = 8'h6F;
Memory[24379] = 8'h6D;
Memory[24378] = 8'h0D;
Memory[24377] = 8'h21;
Memory[24376] = 8'h83;
Memory[24383] = 8'h00;
Memory[24382] = 8'h3B;
Memory[24381] = 8'h2A;
Memory[24380] = 8'h23;
Memory[24387] = 8'h12;
Memory[24386] = 8'h40;
Memory[24385] = 8'h20;
Memory[24384] = 8'h6F;
Memory[24391] = 8'h6D;
Memory[24390] = 8'h4D;
Memory[24389] = 8'h21;
Memory[24388] = 8'h83;
Memory[24395] = 8'h00;
Memory[24394] = 8'h3B;
Memory[24393] = 8'h2A;
Memory[24392] = 8'h23;
Memory[24399] = 8'h12;
Memory[24398] = 8'h40;
Memory[24397] = 8'h20;
Memory[24396] = 8'h6F;
Memory[24403] = 8'h6D;
Memory[24402] = 8'h8D;
Memory[24401] = 8'h21;
Memory[24400] = 8'h83;
Memory[24407] = 8'h00;
Memory[24406] = 8'h3B;
Memory[24405] = 8'h2A;
Memory[24404] = 8'h23;
Memory[24411] = 8'h12;
Memory[24410] = 8'h40;
Memory[24409] = 8'h20;
Memory[24408] = 8'h6F;
Memory[24415] = 8'h6D;
Memory[24414] = 8'hCD;
Memory[24413] = 8'h21;
Memory[24412] = 8'h83;
Memory[24419] = 8'h00;
Memory[24418] = 8'h3B;
Memory[24417] = 8'h2A;
Memory[24416] = 8'h23;
Memory[24423] = 8'h12;
Memory[24422] = 8'h40;
Memory[24421] = 8'h20;
Memory[24420] = 8'h6F;
Memory[24427] = 8'h6E;
Memory[24426] = 8'h0D;
Memory[24425] = 8'h21;
Memory[24424] = 8'h83;
Memory[24431] = 8'h00;
Memory[24430] = 8'h3B;
Memory[24429] = 8'h2A;
Memory[24428] = 8'h23;
Memory[24435] = 8'h12;
Memory[24434] = 8'h40;
Memory[24433] = 8'h20;
Memory[24432] = 8'h6F;
Memory[24439] = 8'h6E;
Memory[24438] = 8'h4D;
Memory[24437] = 8'h21;
Memory[24436] = 8'h83;
Memory[24443] = 8'h00;
Memory[24442] = 8'h3B;
Memory[24441] = 8'h2A;
Memory[24440] = 8'h23;
Memory[24447] = 8'h12;
Memory[24446] = 8'h40;
Memory[24445] = 8'h20;
Memory[24444] = 8'h6F;
Memory[24451] = 8'h03;
Memory[24450] = 8'h40;
Memory[24449] = 8'h01;
Memory[24448] = 8'h13;
Memory[24455] = 8'h00;
Memory[24454] = 8'h0E;
Memory[24453] = 8'h8E;
Memory[24452] = 8'h13;
Memory[24459] = 8'h50;
Memory[24458] = 8'h90;
Memory[24457] = 8'h10;
Memory[24456] = 8'h6F;
Memory[24463] = 8'h00;
Memory[24462] = 8'h00;
Memory[24461] = 8'h00;
Memory[24460] = 8'h00;
Memory[24467] = 8'h00;
Memory[24466] = 8'h00;
Memory[24465] = 8'h00;
Memory[24464] = 8'h00;
Memory[24471] = 8'h00;
Memory[24470] = 8'h00;
Memory[24469] = 8'h00;
Memory[24468] = 8'h00;
Memory[24475] = 8'h00;
Memory[24474] = 8'h00;
Memory[24473] = 8'h00;
Memory[24472] = 8'h00;
Memory[24479] = 8'h00;
Memory[24478] = 8'h00;
Memory[24477] = 8'h00;
Memory[24476] = 8'h00;
Memory[24483] = 8'h00;
Memory[24482] = 8'h00;
Memory[24481] = 8'h00;
Memory[24480] = 8'h00;
Memory[24487] = 8'h00;
Memory[24486] = 8'h00;
Memory[24485] = 8'h00;
Memory[24484] = 8'h00;
Memory[24491] = 8'h00;
Memory[24490] = 8'h00;
Memory[24489] = 8'h00;
Memory[24488] = 8'h00;
Memory[24495] = 8'h00;
Memory[24494] = 8'h00;
Memory[24493] = 8'h00;
Memory[24492] = 8'h00;
Memory[24499] = 8'h00;
Memory[24498] = 8'h00;
Memory[24497] = 8'h00;
Memory[24496] = 8'h00;
Memory[24503] = 8'h00;
Memory[24502] = 8'h00;
Memory[24501] = 8'h00;
Memory[24500] = 8'h00;
Memory[24507] = 8'h00;
Memory[24506] = 8'h00;
Memory[24505] = 8'h00;
Memory[24504] = 8'h00;
Memory[24511] = 8'h00;
Memory[24510] = 8'h00;
Memory[24509] = 8'h00;
Memory[24508] = 8'h00;
Memory[24515] = 8'h00;
Memory[24514] = 8'h00;
Memory[24513] = 8'h00;
Memory[24512] = 8'h00;
Memory[24519] = 8'h00;
Memory[24518] = 8'h00;
Memory[24517] = 8'h00;
Memory[24516] = 8'h00;
Memory[24523] = 8'h00;
Memory[24522] = 8'h00;
Memory[24521] = 8'h00;
Memory[24520] = 8'h00;
Memory[24527] = 8'h00;
Memory[24526] = 8'h00;
Memory[24525] = 8'h00;
Memory[24524] = 8'h00;
Memory[24531] = 8'h00;
Memory[24530] = 8'h00;
Memory[24529] = 8'h00;
Memory[24528] = 8'h00;
Memory[24535] = 8'h00;
Memory[24534] = 8'h00;
Memory[24533] = 8'h00;
Memory[24532] = 8'h00;
Memory[24539] = 8'h00;
Memory[24538] = 8'h00;
Memory[24537] = 8'h00;
Memory[24536] = 8'h00;
Memory[24543] = 8'h00;
Memory[24542] = 8'h00;
Memory[24541] = 8'h00;
Memory[24540] = 8'h00;
Memory[24547] = 8'h00;
Memory[24546] = 8'h00;
Memory[24545] = 8'h00;
Memory[24544] = 8'h00;
Memory[24551] = 8'h00;
Memory[24550] = 8'h00;
Memory[24549] = 8'h00;
Memory[24548] = 8'h00;
Memory[24555] = 8'h00;
Memory[24554] = 8'h00;
Memory[24553] = 8'h00;
Memory[24552] = 8'h00;
Memory[24559] = 8'h00;
Memory[24558] = 8'h00;
Memory[24557] = 8'h00;
Memory[24556] = 8'h00;
Memory[24563] = 8'h00;
Memory[24562] = 8'h00;
Memory[24561] = 8'h00;
Memory[24560] = 8'h00;
Memory[24567] = 8'h00;
Memory[24566] = 8'h00;
Memory[24565] = 8'h00;
Memory[24564] = 8'h00;
Memory[24571] = 8'h00;
Memory[24570] = 8'h00;
Memory[24569] = 8'h00;
Memory[24568] = 8'h00;
Memory[24575] = 8'h00;
Memory[24574] = 8'h00;
Memory[24573] = 8'h00;
Memory[24572] = 8'h00;
Memory[24579] = 8'h00;
Memory[24578] = 8'h00;
Memory[24577] = 8'h00;
Memory[24576] = 8'h00;
Memory[24583] = 8'h00;
Memory[24582] = 8'h00;
Memory[24581] = 8'h00;
Memory[24580] = 8'h00;
Memory[24587] = 8'h00;
Memory[24586] = 8'h00;
Memory[24585] = 8'h00;
Memory[24584] = 8'h00;
Memory[24591] = 8'h00;
Memory[24590] = 8'h00;
Memory[24589] = 8'h00;
Memory[24588] = 8'h00;
Memory[24595] = 8'h00;
Memory[24594] = 8'h00;
Memory[24593] = 8'h00;
Memory[24592] = 8'h00;
Memory[24599] = 8'h00;
Memory[24598] = 8'h00;
Memory[24597] = 8'h00;
Memory[24596] = 8'h00;
Memory[24603] = 8'h00;
Memory[24602] = 8'h00;
Memory[24601] = 8'h00;
Memory[24600] = 8'h00;
Memory[24607] = 8'h00;
Memory[24606] = 8'h00;
Memory[24605] = 8'h00;
Memory[24604] = 8'h00;
Memory[24611] = 8'h00;
Memory[24610] = 8'h00;
Memory[24609] = 8'h00;
Memory[24608] = 8'h00;
Memory[24615] = 8'h00;
Memory[24614] = 8'h00;
Memory[24613] = 8'h00;
Memory[24612] = 8'h00;
Memory[24619] = 8'h00;
Memory[24618] = 8'h00;
Memory[24617] = 8'h00;
Memory[24616] = 8'h00;
Memory[24623] = 8'h00;
Memory[24622] = 8'h00;
Memory[24621] = 8'h00;
Memory[24620] = 8'h00;
Memory[24627] = 8'h00;
Memory[24626] = 8'h00;
Memory[24625] = 8'h00;
Memory[24624] = 8'h00;
Memory[24631] = 8'h00;
Memory[24630] = 8'h00;
Memory[24629] = 8'h00;
Memory[24628] = 8'h00;
Memory[24635] = 8'h00;
Memory[24634] = 8'h00;
Memory[24633] = 8'h00;
Memory[24632] = 8'h00;
Memory[24639] = 8'h00;
Memory[24638] = 8'h00;
Memory[24637] = 8'h00;
Memory[24636] = 8'h00;
Memory[24643] = 8'h00;
Memory[24642] = 8'h00;
Memory[24641] = 8'h00;
Memory[24640] = 8'h00;
Memory[24647] = 8'h00;
Memory[24646] = 8'h00;
Memory[24645] = 8'h00;
Memory[24644] = 8'h00;
Memory[24651] = 8'h00;
Memory[24650] = 8'h00;
Memory[24649] = 8'h00;
Memory[24648] = 8'h00;
Memory[24655] = 8'h00;
Memory[24654] = 8'h00;
Memory[24653] = 8'h00;
Memory[24652] = 8'h00;
Memory[24659] = 8'h00;
Memory[24658] = 8'h00;
Memory[24657] = 8'h00;
Memory[24656] = 8'h00;
Memory[24663] = 8'h00;
Memory[24662] = 8'h00;
Memory[24661] = 8'h00;
Memory[24660] = 8'h00;
Memory[24667] = 8'h00;
Memory[24666] = 8'h00;
Memory[24665] = 8'h00;
Memory[24664] = 8'h00;
Memory[24671] = 8'h00;
Memory[24670] = 8'h00;
Memory[24669] = 8'h00;
Memory[24668] = 8'h00;
Memory[24675] = 8'h00;
Memory[24674] = 8'h00;
Memory[24673] = 8'h00;
Memory[24672] = 8'h00;
Memory[24679] = 8'h00;
Memory[24678] = 8'h00;
Memory[24677] = 8'h00;
Memory[24676] = 8'h00;
Memory[24683] = 8'h00;
Memory[24682] = 8'h00;
Memory[24681] = 8'h00;
Memory[24680] = 8'h00;
Memory[24687] = 8'h00;
Memory[24686] = 8'h00;
Memory[24685] = 8'h00;
Memory[24684] = 8'h00;
Memory[24691] = 8'h00;
Memory[24690] = 8'h00;
Memory[24689] = 8'h00;
Memory[24688] = 8'h00;
Memory[24695] = 8'h00;
Memory[24694] = 8'h00;
Memory[24693] = 8'h00;
Memory[24692] = 8'h00;
Memory[24699] = 8'h00;
Memory[24698] = 8'h00;
Memory[24697] = 8'h00;
Memory[24696] = 8'h00;
Memory[24703] = 8'h00;
Memory[24702] = 8'h00;
Memory[24701] = 8'h00;
Memory[24700] = 8'h00;
Memory[24707] = 8'h00;
Memory[24706] = 8'h00;
Memory[24705] = 8'h00;
Memory[24704] = 8'h00;
Memory[24711] = 8'h00;
Memory[24710] = 8'h00;
Memory[24709] = 8'h00;
Memory[24708] = 8'h00;
Memory[24715] = 8'h00;
Memory[24714] = 8'h00;
Memory[24713] = 8'h00;
Memory[24712] = 8'h00;
Memory[24719] = 8'h00;
Memory[24718] = 8'h00;
Memory[24717] = 8'h00;
Memory[24716] = 8'h00;
Memory[24723] = 8'h00;
Memory[24722] = 8'h00;
Memory[24721] = 8'h00;
Memory[24720] = 8'h00;
Memory[24727] = 8'h00;
Memory[24726] = 8'h00;
Memory[24725] = 8'h00;
Memory[24724] = 8'h00;
Memory[24731] = 8'h00;
Memory[24730] = 8'h00;
Memory[24729] = 8'h00;
Memory[24728] = 8'h00;
Memory[24735] = 8'h00;
Memory[24734] = 8'h00;
Memory[24733] = 8'h00;
Memory[24732] = 8'h00;
Memory[24739] = 8'h00;
Memory[24738] = 8'h00;
Memory[24737] = 8'h00;
Memory[24736] = 8'h00;
Memory[24743] = 8'h00;
Memory[24742] = 8'h00;
Memory[24741] = 8'h00;
Memory[24740] = 8'h00;
Memory[24747] = 8'h00;
Memory[24746] = 8'h00;
Memory[24745] = 8'h00;
Memory[24744] = 8'h00;
Memory[24751] = 8'h00;
Memory[24750] = 8'h00;
Memory[24749] = 8'h00;
Memory[24748] = 8'h00;
Memory[24755] = 8'h00;
Memory[24754] = 8'h00;
Memory[24753] = 8'h00;
Memory[24752] = 8'h00;
Memory[24759] = 8'h00;
Memory[24758] = 8'h00;
Memory[24757] = 8'h00;
Memory[24756] = 8'h00;
Memory[24763] = 8'h00;
Memory[24762] = 8'h00;
Memory[24761] = 8'h00;
Memory[24760] = 8'h00;
Memory[24767] = 8'h00;
Memory[24766] = 8'h00;
Memory[24765] = 8'h00;
Memory[24764] = 8'h00;
Memory[24771] = 8'h00;
Memory[24770] = 8'h00;
Memory[24769] = 8'h00;
Memory[24768] = 8'h00;
Memory[24775] = 8'h00;
Memory[24774] = 8'h00;
Memory[24773] = 8'h00;
Memory[24772] = 8'h00;
Memory[24779] = 8'h00;
Memory[24778] = 8'h00;
Memory[24777] = 8'h00;
Memory[24776] = 8'h00;
Memory[24783] = 8'h00;
Memory[24782] = 8'h00;
Memory[24781] = 8'h00;
Memory[24780] = 8'h00;
Memory[24787] = 8'h00;
Memory[24786] = 8'h00;
Memory[24785] = 8'h00;
Memory[24784] = 8'h00;
Memory[24791] = 8'h00;
Memory[24790] = 8'h00;
Memory[24789] = 8'h00;
Memory[24788] = 8'h00;
Memory[24795] = 8'h00;
Memory[24794] = 8'h00;
Memory[24793] = 8'h00;
Memory[24792] = 8'h00;
Memory[24799] = 8'h00;
Memory[24798] = 8'h00;
Memory[24797] = 8'h00;
Memory[24796] = 8'h00;
Memory[24803] = 8'h00;
Memory[24802] = 8'h00;
Memory[24801] = 8'h00;
Memory[24800] = 8'h00;
Memory[24807] = 8'h00;
Memory[24806] = 8'h00;
Memory[24805] = 8'h00;
Memory[24804] = 8'h00;
Memory[24811] = 8'h00;
Memory[24810] = 8'h00;
Memory[24809] = 8'h00;
Memory[24808] = 8'h00;
Memory[24815] = 8'h00;
Memory[24814] = 8'h00;
Memory[24813] = 8'h00;
Memory[24812] = 8'h00;
Memory[24819] = 8'h00;
Memory[24818] = 8'h00;
Memory[24817] = 8'h00;
Memory[24816] = 8'h00;
Memory[24823] = 8'h00;
Memory[24822] = 8'h00;
Memory[24821] = 8'h00;
Memory[24820] = 8'h00;
Memory[24827] = 8'h00;
Memory[24826] = 8'h00;
Memory[24825] = 8'h00;
Memory[24824] = 8'h00;
Memory[24831] = 8'h00;
Memory[24830] = 8'h00;
Memory[24829] = 8'h00;
Memory[24828] = 8'h00;
Memory[24835] = 8'h00;
Memory[24834] = 8'h00;
Memory[24833] = 8'h00;
Memory[24832] = 8'h00;
Memory[24839] = 8'h00;
Memory[24838] = 8'h00;
Memory[24837] = 8'h00;
Memory[24836] = 8'h00;
Memory[24843] = 8'h00;
Memory[24842] = 8'h00;
Memory[24841] = 8'h00;
Memory[24840] = 8'h00;
Memory[24847] = 8'h00;
Memory[24846] = 8'h00;
Memory[24845] = 8'h00;
Memory[24844] = 8'h00;
Memory[24851] = 8'h00;
Memory[24850] = 8'h00;
Memory[24849] = 8'h00;
Memory[24848] = 8'h00;
Memory[24855] = 8'h00;
Memory[24854] = 8'h00;
Memory[24853] = 8'h00;
Memory[24852] = 8'h00;
Memory[24859] = 8'h00;
Memory[24858] = 8'h00;
Memory[24857] = 8'h00;
Memory[24856] = 8'h00;
Memory[24863] = 8'h00;
Memory[24862] = 8'h00;
Memory[24861] = 8'h00;
Memory[24860] = 8'h00;
Memory[24867] = 8'h00;
Memory[24866] = 8'h00;
Memory[24865] = 8'h00;
Memory[24864] = 8'h00;
Memory[24871] = 8'h00;
Memory[24870] = 8'h00;
Memory[24869] = 8'h00;
Memory[24868] = 8'h00;
Memory[24875] = 8'h00;
Memory[24874] = 8'h00;
Memory[24873] = 8'h00;
Memory[24872] = 8'h00;
Memory[24879] = 8'h00;
Memory[24878] = 8'h00;
Memory[24877] = 8'h00;
Memory[24876] = 8'h00;
Memory[24883] = 8'h00;
Memory[24882] = 8'h00;
Memory[24881] = 8'h00;
Memory[24880] = 8'h00;
Memory[24887] = 8'h00;
Memory[24886] = 8'h00;
Memory[24885] = 8'h00;
Memory[24884] = 8'h00;
Memory[24891] = 8'h00;
Memory[24890] = 8'h00;
Memory[24889] = 8'h00;
Memory[24888] = 8'h00;
Memory[24895] = 8'h00;
Memory[24894] = 8'h00;
Memory[24893] = 8'h00;
Memory[24892] = 8'h00;
Memory[24899] = 8'h00;
Memory[24898] = 8'h00;
Memory[24897] = 8'h00;
Memory[24896] = 8'h00;
Memory[24903] = 8'h00;
Memory[24902] = 8'h00;
Memory[24901] = 8'h00;
Memory[24900] = 8'h00;
Memory[24907] = 8'h00;
Memory[24906] = 8'h00;
Memory[24905] = 8'h00;
Memory[24904] = 8'h00;
Memory[24911] = 8'h00;
Memory[24910] = 8'h00;
Memory[24909] = 8'h00;
Memory[24908] = 8'h00;
Memory[24915] = 8'h00;
Memory[24914] = 8'h00;
Memory[24913] = 8'h00;
Memory[24912] = 8'h00;
Memory[24919] = 8'h00;
Memory[24918] = 8'h00;
Memory[24917] = 8'h00;
Memory[24916] = 8'h00;
Memory[24923] = 8'h00;
Memory[24922] = 8'h00;
Memory[24921] = 8'h00;
Memory[24920] = 8'h00;
Memory[24927] = 8'h00;
Memory[24926] = 8'h00;
Memory[24925] = 8'h00;
Memory[24924] = 8'h00;
Memory[24931] = 8'h00;
Memory[24930] = 8'h00;
Memory[24929] = 8'h00;
Memory[24928] = 8'h00;
Memory[24935] = 8'h00;
Memory[24934] = 8'h00;
Memory[24933] = 8'h00;
Memory[24932] = 8'h00;
Memory[24939] = 8'h00;
Memory[24938] = 8'h00;
Memory[24937] = 8'h00;
Memory[24936] = 8'h00;
Memory[24943] = 8'h00;
Memory[24942] = 8'h00;
Memory[24941] = 8'h00;
Memory[24940] = 8'h00;
Memory[24947] = 8'h00;
Memory[24946] = 8'h00;
Memory[24945] = 8'h00;
Memory[24944] = 8'h00;
Memory[24951] = 8'h00;
Memory[24950] = 8'h00;
Memory[24949] = 8'h00;
Memory[24948] = 8'h00;
Memory[24955] = 8'h00;
Memory[24954] = 8'h00;
Memory[24953] = 8'h00;
Memory[24952] = 8'h00;
Memory[24959] = 8'h00;
Memory[24958] = 8'h00;
Memory[24957] = 8'h00;
Memory[24956] = 8'h00;
Memory[24963] = 8'h00;
Memory[24962] = 8'h00;
Memory[24961] = 8'h00;
Memory[24960] = 8'h00;
Memory[24967] = 8'h00;
Memory[24966] = 8'h00;
Memory[24965] = 8'h00;
Memory[24964] = 8'h00;
Memory[24971] = 8'h00;
Memory[24970] = 8'h00;
Memory[24969] = 8'h00;
Memory[24968] = 8'h00;
Memory[24975] = 8'h00;
Memory[24974] = 8'h00;
Memory[24973] = 8'h00;
Memory[24972] = 8'h00;
Memory[24979] = 8'h00;
Memory[24978] = 8'h00;
Memory[24977] = 8'h00;
Memory[24976] = 8'h00;
Memory[24983] = 8'h00;
Memory[24982] = 8'h00;
Memory[24981] = 8'h00;
Memory[24980] = 8'h00;
Memory[24987] = 8'h00;
Memory[24986] = 8'h00;
Memory[24985] = 8'h00;
Memory[24984] = 8'h00;
Memory[24991] = 8'h00;
Memory[24990] = 8'h00;
Memory[24989] = 8'h00;
Memory[24988] = 8'h00;
Memory[24995] = 8'h00;
Memory[24994] = 8'h00;
Memory[24993] = 8'h00;
Memory[24992] = 8'h00;
Memory[24999] = 8'h00;
Memory[24998] = 8'h00;
Memory[24997] = 8'h00;
Memory[24996] = 8'h00;
Memory[25003] = 8'h00;
Memory[25002] = 8'h00;
Memory[25001] = 8'h00;
Memory[25000] = 8'h00;
Memory[25007] = 8'h00;
Memory[25006] = 8'h00;
Memory[25005] = 8'h00;
Memory[25004] = 8'h00;
Memory[25011] = 8'h00;
Memory[25010] = 8'h00;
Memory[25009] = 8'h00;
Memory[25008] = 8'h00;
Memory[25015] = 8'h00;
Memory[25014] = 8'h00;
Memory[25013] = 8'h00;
Memory[25012] = 8'h00;
Memory[25019] = 8'h00;
Memory[25018] = 8'h00;
Memory[25017] = 8'h00;
Memory[25016] = 8'h00;
Memory[25023] = 8'h00;
Memory[25022] = 8'h00;
Memory[25021] = 8'h00;
Memory[25020] = 8'h00;
Memory[25027] = 8'h00;
Memory[25026] = 8'h00;
Memory[25025] = 8'h00;
Memory[25024] = 8'h00;
Memory[25031] = 8'h00;
Memory[25030] = 8'h00;
Memory[25029] = 8'h00;
Memory[25028] = 8'h00;
Memory[25035] = 8'h00;
Memory[25034] = 8'h00;
Memory[25033] = 8'h00;
Memory[25032] = 8'h00;
Memory[25039] = 8'h00;
Memory[25038] = 8'h00;
Memory[25037] = 8'h00;
Memory[25036] = 8'h00;
Memory[25043] = 8'h00;
Memory[25042] = 8'h00;
Memory[25041] = 8'h00;
Memory[25040] = 8'h00;
Memory[25047] = 8'h00;
Memory[25046] = 8'h00;
Memory[25045] = 8'h00;
Memory[25044] = 8'h00;
Memory[25051] = 8'h00;
Memory[25050] = 8'h00;
Memory[25049] = 8'h00;
Memory[25048] = 8'h00;
Memory[25055] = 8'h00;
Memory[25054] = 8'h00;
Memory[25053] = 8'h00;
Memory[25052] = 8'h00;
Memory[25059] = 8'h00;
Memory[25058] = 8'h00;
Memory[25057] = 8'h00;
Memory[25056] = 8'h00;
Memory[25063] = 8'h00;
Memory[25062] = 8'h00;
Memory[25061] = 8'h00;
Memory[25060] = 8'h00;
Memory[25067] = 8'h00;
Memory[25066] = 8'h00;
Memory[25065] = 8'h00;
Memory[25064] = 8'h00;
Memory[25071] = 8'h00;
Memory[25070] = 8'h00;
Memory[25069] = 8'h00;
Memory[25068] = 8'h00;
Memory[25075] = 8'h00;
Memory[25074] = 8'h00;
Memory[25073] = 8'h00;
Memory[25072] = 8'h00;
Memory[25079] = 8'h00;
Memory[25078] = 8'h00;
Memory[25077] = 8'h00;
Memory[25076] = 8'h00;
Memory[25083] = 8'h00;
Memory[25082] = 8'h00;
Memory[25081] = 8'h00;
Memory[25080] = 8'h00;
Memory[25087] = 8'h00;
Memory[25086] = 8'h00;
Memory[25085] = 8'h00;
Memory[25084] = 8'h00;
Memory[25091] = 8'h00;
Memory[25090] = 8'h00;
Memory[25089] = 8'h00;
Memory[25088] = 8'h00;
Memory[25095] = 8'h00;
Memory[25094] = 8'h00;
Memory[25093] = 8'h00;
Memory[25092] = 8'h00;
Memory[25099] = 8'h00;
Memory[25098] = 8'h00;
Memory[25097] = 8'h00;
Memory[25096] = 8'h00;
Memory[25103] = 8'h00;
Memory[25102] = 8'h00;
Memory[25101] = 8'h00;
Memory[25100] = 8'h00;
Memory[25107] = 8'h00;
Memory[25106] = 8'h00;
Memory[25105] = 8'h00;
Memory[25104] = 8'h00;
Memory[25111] = 8'h00;
Memory[25110] = 8'h00;
Memory[25109] = 8'h00;
Memory[25108] = 8'h00;
Memory[25115] = 8'h00;
Memory[25114] = 8'h00;
Memory[25113] = 8'h00;
Memory[25112] = 8'h00;
Memory[25119] = 8'h00;
Memory[25118] = 8'h00;
Memory[25117] = 8'h00;
Memory[25116] = 8'h00;
Memory[25123] = 8'h00;
Memory[25122] = 8'h00;
Memory[25121] = 8'h00;
Memory[25120] = 8'h00;
Memory[25127] = 8'h00;
Memory[25126] = 8'h00;
Memory[25125] = 8'h00;
Memory[25124] = 8'h00;
Memory[25131] = 8'h00;
Memory[25130] = 8'h00;
Memory[25129] = 8'h00;
Memory[25128] = 8'h00;
Memory[25135] = 8'h00;
Memory[25134] = 8'h00;
Memory[25133] = 8'h00;
Memory[25132] = 8'h00;
Memory[25139] = 8'h00;
Memory[25138] = 8'h00;
Memory[25137] = 8'h00;
Memory[25136] = 8'h00;
Memory[25143] = 8'h00;
Memory[25142] = 8'h00;
Memory[25141] = 8'h00;
Memory[25140] = 8'h00;
Memory[25147] = 8'h00;
Memory[25146] = 8'h00;
Memory[25145] = 8'h00;
Memory[25144] = 8'h00;
Memory[25151] = 8'h00;
Memory[25150] = 8'h00;
Memory[25149] = 8'h00;
Memory[25148] = 8'h00;
Memory[25155] = 8'h00;
Memory[25154] = 8'h00;
Memory[25153] = 8'h00;
Memory[25152] = 8'h00;
Memory[25159] = 8'h00;
Memory[25158] = 8'h00;
Memory[25157] = 8'h00;
Memory[25156] = 8'h00;
Memory[25163] = 8'h00;
Memory[25162] = 8'h00;
Memory[25161] = 8'h00;
Memory[25160] = 8'h00;
Memory[25167] = 8'h00;
Memory[25166] = 8'h00;
Memory[25165] = 8'h00;
Memory[25164] = 8'h00;
Memory[25171] = 8'h00;
Memory[25170] = 8'h00;
Memory[25169] = 8'h00;
Memory[25168] = 8'h00;
Memory[25175] = 8'h00;
Memory[25174] = 8'h00;
Memory[25173] = 8'h00;
Memory[25172] = 8'h00;
Memory[25179] = 8'h00;
Memory[25178] = 8'h00;
Memory[25177] = 8'h00;
Memory[25176] = 8'h00;
Memory[25183] = 8'h00;
Memory[25182] = 8'h00;
Memory[25181] = 8'h00;
Memory[25180] = 8'h00;
Memory[25187] = 8'h00;
Memory[25186] = 8'h00;
Memory[25185] = 8'h00;
Memory[25184] = 8'h00;
Memory[25191] = 8'h00;
Memory[25190] = 8'h00;
Memory[25189] = 8'h00;
Memory[25188] = 8'h00;
Memory[25195] = 8'h00;
Memory[25194] = 8'h00;
Memory[25193] = 8'h00;
Memory[25192] = 8'h00;
Memory[25199] = 8'h00;
Memory[25198] = 8'h00;
Memory[25197] = 8'h00;
Memory[25196] = 8'h00;
Memory[25203] = 8'h00;
Memory[25202] = 8'h00;
Memory[25201] = 8'h00;
Memory[25200] = 8'h00;
Memory[25207] = 8'h00;
Memory[25206] = 8'h00;
Memory[25205] = 8'h00;
Memory[25204] = 8'h00;
Memory[25211] = 8'h00;
Memory[25210] = 8'h00;
Memory[25209] = 8'h00;
Memory[25208] = 8'h00;
Memory[25215] = 8'h00;
Memory[25214] = 8'h00;
Memory[25213] = 8'h00;
Memory[25212] = 8'h00;
Memory[25219] = 8'h00;
Memory[25218] = 8'h00;
Memory[25217] = 8'h00;
Memory[25216] = 8'h00;
Memory[25223] = 8'h00;
Memory[25222] = 8'h00;
Memory[25221] = 8'h00;
Memory[25220] = 8'h00;
Memory[25227] = 8'h00;
Memory[25226] = 8'h00;
Memory[25225] = 8'h00;
Memory[25224] = 8'h00;
Memory[25231] = 8'h00;
Memory[25230] = 8'h00;
Memory[25229] = 8'h00;
Memory[25228] = 8'h00;
Memory[25235] = 8'h00;
Memory[25234] = 8'h00;
Memory[25233] = 8'h00;
Memory[25232] = 8'h00;
Memory[25239] = 8'h00;
Memory[25238] = 8'h00;
Memory[25237] = 8'h00;
Memory[25236] = 8'h00;
Memory[25243] = 8'h00;
Memory[25242] = 8'h00;
Memory[25241] = 8'h00;
Memory[25240] = 8'h00;
Memory[25247] = 8'h00;
Memory[25246] = 8'h00;
Memory[25245] = 8'h00;
Memory[25244] = 8'h00;
Memory[25251] = 8'h00;
Memory[25250] = 8'h00;
Memory[25249] = 8'h00;
Memory[25248] = 8'h00;
Memory[25255] = 8'h00;
Memory[25254] = 8'h00;
Memory[25253] = 8'h00;
Memory[25252] = 8'h00;
Memory[25259] = 8'h00;
Memory[25258] = 8'h00;
Memory[25257] = 8'h00;
Memory[25256] = 8'h00;
Memory[25263] = 8'h00;
Memory[25262] = 8'h00;
Memory[25261] = 8'h00;
Memory[25260] = 8'h00;
Memory[25267] = 8'h00;
Memory[25266] = 8'h00;
Memory[25265] = 8'h00;
Memory[25264] = 8'h00;
Memory[25271] = 8'h00;
Memory[25270] = 8'h00;
Memory[25269] = 8'h00;
Memory[25268] = 8'h00;
Memory[25275] = 8'h00;
Memory[25274] = 8'h00;
Memory[25273] = 8'h00;
Memory[25272] = 8'h00;
Memory[25279] = 8'h00;
Memory[25278] = 8'h00;
Memory[25277] = 8'h00;
Memory[25276] = 8'h00;
Memory[25283] = 8'h00;
Memory[25282] = 8'h00;
Memory[25281] = 8'h00;
Memory[25280] = 8'h00;
Memory[25287] = 8'h00;
Memory[25286] = 8'h00;
Memory[25285] = 8'h00;
Memory[25284] = 8'h00;
Memory[25291] = 8'h00;
Memory[25290] = 8'h00;
Memory[25289] = 8'h00;
Memory[25288] = 8'h00;
Memory[25295] = 8'h00;
Memory[25294] = 8'h00;
Memory[25293] = 8'h00;
Memory[25292] = 8'h00;
Memory[25299] = 8'h00;
Memory[25298] = 8'h00;
Memory[25297] = 8'h00;
Memory[25296] = 8'h00;
Memory[25303] = 8'h00;
Memory[25302] = 8'h00;
Memory[25301] = 8'h00;
Memory[25300] = 8'h00;
Memory[25307] = 8'h00;
Memory[25306] = 8'h00;
Memory[25305] = 8'h00;
Memory[25304] = 8'h00;
Memory[25311] = 8'h00;
Memory[25310] = 8'h00;
Memory[25309] = 8'h00;
Memory[25308] = 8'h00;
Memory[25315] = 8'h00;
Memory[25314] = 8'h00;
Memory[25313] = 8'h00;
Memory[25312] = 8'h00;
Memory[25319] = 8'h00;
Memory[25318] = 8'h00;
Memory[25317] = 8'h00;
Memory[25316] = 8'h00;
Memory[25323] = 8'h00;
Memory[25322] = 8'h00;
Memory[25321] = 8'h00;
Memory[25320] = 8'h00;
Memory[25327] = 8'h00;
Memory[25326] = 8'h00;
Memory[25325] = 8'h00;
Memory[25324] = 8'h00;
Memory[25331] = 8'h00;
Memory[25330] = 8'h00;
Memory[25329] = 8'h00;
Memory[25328] = 8'h00;
Memory[25335] = 8'h00;
Memory[25334] = 8'h00;
Memory[25333] = 8'h00;
Memory[25332] = 8'h00;
Memory[25339] = 8'h00;
Memory[25338] = 8'h00;
Memory[25337] = 8'h00;
Memory[25336] = 8'h00;
Memory[25343] = 8'h00;
Memory[25342] = 8'h00;
Memory[25341] = 8'h00;
Memory[25340] = 8'h00;
Memory[25347] = 8'h00;
Memory[25346] = 8'h00;
Memory[25345] = 8'h00;
Memory[25344] = 8'h00;
Memory[25351] = 8'h00;
Memory[25350] = 8'h00;
Memory[25349] = 8'h00;
Memory[25348] = 8'h00;
Memory[25355] = 8'h00;
Memory[25354] = 8'h00;
Memory[25353] = 8'h00;
Memory[25352] = 8'h00;
Memory[25359] = 8'h00;
Memory[25358] = 8'h00;
Memory[25357] = 8'h00;
Memory[25356] = 8'h00;
Memory[25363] = 8'h00;
Memory[25362] = 8'h00;
Memory[25361] = 8'h00;
Memory[25360] = 8'h00;
Memory[25367] = 8'h00;
Memory[25366] = 8'h00;
Memory[25365] = 8'h00;
Memory[25364] = 8'h00;
Memory[25371] = 8'h00;
Memory[25370] = 8'h00;
Memory[25369] = 8'h00;
Memory[25368] = 8'h00;
Memory[25375] = 8'h00;
Memory[25374] = 8'h00;
Memory[25373] = 8'h00;
Memory[25372] = 8'h00;
Memory[25379] = 8'h00;
Memory[25378] = 8'h00;
Memory[25377] = 8'h00;
Memory[25376] = 8'h00;
Memory[25383] = 8'h00;
Memory[25382] = 8'h00;
Memory[25381] = 8'h00;
Memory[25380] = 8'h00;
Memory[25387] = 8'h00;
Memory[25386] = 8'h00;
Memory[25385] = 8'h00;
Memory[25384] = 8'h00;
Memory[25391] = 8'h00;
Memory[25390] = 8'h00;
Memory[25389] = 8'h00;
Memory[25388] = 8'h00;
Memory[25395] = 8'h00;
Memory[25394] = 8'h00;
Memory[25393] = 8'h00;
Memory[25392] = 8'h00;
Memory[25399] = 8'h00;
Memory[25398] = 8'h00;
Memory[25397] = 8'h00;
Memory[25396] = 8'h00;
Memory[25403] = 8'h00;
Memory[25402] = 8'h00;
Memory[25401] = 8'h00;
Memory[25400] = 8'h00;
Memory[25407] = 8'h00;
Memory[25406] = 8'h00;
Memory[25405] = 8'h00;
Memory[25404] = 8'h00;
Memory[25411] = 8'h00;
Memory[25410] = 8'h00;
Memory[25409] = 8'h00;
Memory[25408] = 8'h00;
Memory[25415] = 8'h00;
Memory[25414] = 8'h00;
Memory[25413] = 8'h00;
Memory[25412] = 8'h00;
Memory[25419] = 8'h00;
Memory[25418] = 8'h00;
Memory[25417] = 8'h00;
Memory[25416] = 8'h00;
Memory[25423] = 8'h00;
Memory[25422] = 8'h00;
Memory[25421] = 8'h00;
Memory[25420] = 8'h00;
Memory[25427] = 8'h00;
Memory[25426] = 8'h00;
Memory[25425] = 8'h00;
Memory[25424] = 8'h00;
Memory[25431] = 8'h00;
Memory[25430] = 8'h00;
Memory[25429] = 8'h00;
Memory[25428] = 8'h00;
Memory[25435] = 8'h00;
Memory[25434] = 8'h00;
Memory[25433] = 8'h00;
Memory[25432] = 8'h00;
Memory[25439] = 8'h00;
Memory[25438] = 8'h00;
Memory[25437] = 8'h00;
Memory[25436] = 8'h00;
Memory[25443] = 8'h00;
Memory[25442] = 8'h00;
Memory[25441] = 8'h00;
Memory[25440] = 8'h00;
Memory[25447] = 8'h00;
Memory[25446] = 8'h00;
Memory[25445] = 8'h00;
Memory[25444] = 8'h00;
Memory[25451] = 8'h00;
Memory[25450] = 8'h00;
Memory[25449] = 8'h00;
Memory[25448] = 8'h00;
Memory[25455] = 8'h00;
Memory[25454] = 8'h00;
Memory[25453] = 8'h00;
Memory[25452] = 8'h00;
Memory[25459] = 8'h00;
Memory[25458] = 8'h00;
Memory[25457] = 8'h00;
Memory[25456] = 8'h00;
Memory[25463] = 8'h00;
Memory[25462] = 8'h00;
Memory[25461] = 8'h00;
Memory[25460] = 8'h00;
Memory[25467] = 8'h00;
Memory[25466] = 8'h00;
Memory[25465] = 8'h00;
Memory[25464] = 8'h00;
Memory[25471] = 8'h00;
Memory[25470] = 8'h00;
Memory[25469] = 8'h00;
Memory[25468] = 8'h00;
Memory[25475] = 8'h00;
Memory[25474] = 8'h00;
Memory[25473] = 8'h00;
Memory[25472] = 8'h00;
Memory[25479] = 8'h00;
Memory[25478] = 8'h00;
Memory[25477] = 8'h00;
Memory[25476] = 8'h00;
Memory[25483] = 8'h00;
Memory[25482] = 8'h00;
Memory[25481] = 8'h00;
Memory[25480] = 8'h00;
Memory[25487] = 8'h00;
Memory[25486] = 8'h00;
Memory[25485] = 8'h00;
Memory[25484] = 8'h00;
Memory[25491] = 8'h00;
Memory[25490] = 8'h00;
Memory[25489] = 8'h00;
Memory[25488] = 8'h00;
Memory[25495] = 8'h00;
Memory[25494] = 8'h00;
Memory[25493] = 8'h00;
Memory[25492] = 8'h00;
Memory[25499] = 8'h00;
Memory[25498] = 8'h00;
Memory[25497] = 8'h00;
Memory[25496] = 8'h00;
Memory[25503] = 8'h00;
Memory[25502] = 8'h00;
Memory[25501] = 8'h00;
Memory[25500] = 8'h00;
Memory[25507] = 8'h00;
Memory[25506] = 8'h00;
Memory[25505] = 8'h00;
Memory[25504] = 8'h00;
Memory[25511] = 8'h00;
Memory[25510] = 8'h00;
Memory[25509] = 8'h00;
Memory[25508] = 8'h00;
Memory[25515] = 8'h00;
Memory[25514] = 8'h00;
Memory[25513] = 8'h00;
Memory[25512] = 8'h00;
Memory[25519] = 8'h00;
Memory[25518] = 8'h00;
Memory[25517] = 8'h00;
Memory[25516] = 8'h00;
Memory[25523] = 8'h00;
Memory[25522] = 8'h00;
Memory[25521] = 8'h00;
Memory[25520] = 8'h00;
Memory[25527] = 8'h00;
Memory[25526] = 8'h00;
Memory[25525] = 8'h00;
Memory[25524] = 8'h00;
Memory[25531] = 8'h00;
Memory[25530] = 8'h00;
Memory[25529] = 8'h00;
Memory[25528] = 8'h00;
Memory[25535] = 8'h00;
Memory[25534] = 8'h00;
Memory[25533] = 8'h00;
Memory[25532] = 8'h00;
Memory[25539] = 8'h00;
Memory[25538] = 8'h00;
Memory[25537] = 8'h00;
Memory[25536] = 8'h00;
Memory[25543] = 8'h00;
Memory[25542] = 8'h00;
Memory[25541] = 8'h00;
Memory[25540] = 8'h00;
Memory[25547] = 8'h00;
Memory[25546] = 8'h00;
Memory[25545] = 8'h00;
Memory[25544] = 8'h00;
Memory[25551] = 8'h00;
Memory[25550] = 8'h00;
Memory[25549] = 8'h00;
Memory[25548] = 8'h00;
Memory[25555] = 8'h00;
Memory[25554] = 8'h00;
Memory[25553] = 8'h00;
Memory[25552] = 8'h00;
Memory[25559] = 8'h00;
Memory[25558] = 8'h00;
Memory[25557] = 8'h00;
Memory[25556] = 8'h00;
Memory[25563] = 8'h00;
Memory[25562] = 8'h00;
Memory[25561] = 8'h00;
Memory[25560] = 8'h00;
Memory[25567] = 8'h00;
Memory[25566] = 8'h00;
Memory[25565] = 8'h00;
Memory[25564] = 8'h00;
Memory[25571] = 8'h00;
Memory[25570] = 8'h00;
Memory[25569] = 8'h00;
Memory[25568] = 8'h00;
Memory[25575] = 8'h00;
Memory[25574] = 8'h00;
Memory[25573] = 8'h00;
Memory[25572] = 8'h00;
Memory[25579] = 8'h00;
Memory[25578] = 8'h00;
Memory[25577] = 8'h00;
Memory[25576] = 8'h00;
Memory[25583] = 8'h00;
Memory[25582] = 8'h00;
Memory[25581] = 8'h00;
Memory[25580] = 8'h00;
Memory[25587] = 8'h00;
Memory[25586] = 8'h00;
Memory[25585] = 8'h00;
Memory[25584] = 8'h00;
Memory[25591] = 8'h00;
Memory[25590] = 8'h00;
Memory[25589] = 8'h00;
Memory[25588] = 8'h00;
Memory[25595] = 8'h00;
Memory[25594] = 8'h00;
Memory[25593] = 8'h00;
Memory[25592] = 8'h00;
Memory[25599] = 8'h00;
Memory[25598] = 8'h00;
Memory[25597] = 8'h00;
Memory[25596] = 8'h00;
Memory[25603] = 8'h00;
Memory[25602] = 8'h00;
Memory[25601] = 8'h00;
Memory[25600] = 8'h00;
Memory[25607] = 8'h00;
Memory[25606] = 8'h00;
Memory[25605] = 8'h00;
Memory[25604] = 8'h00;
Memory[25611] = 8'h00;
Memory[25610] = 8'h00;
Memory[25609] = 8'h00;
Memory[25608] = 8'h00;
Memory[25615] = 8'h00;
Memory[25614] = 8'h00;
Memory[25613] = 8'h00;
Memory[25612] = 8'h00;
Memory[25619] = 8'h00;
Memory[25618] = 8'h00;
Memory[25617] = 8'h00;
Memory[25616] = 8'h00;
Memory[25623] = 8'h00;
Memory[25622] = 8'h00;
Memory[25621] = 8'h00;
Memory[25620] = 8'h00;
Memory[25627] = 8'h00;
Memory[25626] = 8'h00;
Memory[25625] = 8'h00;
Memory[25624] = 8'h00;
Memory[25631] = 8'h00;
Memory[25630] = 8'h00;
Memory[25629] = 8'h00;
Memory[25628] = 8'h00;
Memory[25635] = 8'h00;
Memory[25634] = 8'h00;
Memory[25633] = 8'h00;
Memory[25632] = 8'h00;
Memory[25639] = 8'h00;
Memory[25638] = 8'h00;
Memory[25637] = 8'h00;
Memory[25636] = 8'h00;
Memory[25643] = 8'h00;
Memory[25642] = 8'h00;
Memory[25641] = 8'h00;
Memory[25640] = 8'h00;
Memory[25647] = 8'h00;
Memory[25646] = 8'h00;
Memory[25645] = 8'h00;
Memory[25644] = 8'h00;
Memory[25651] = 8'h00;
Memory[25650] = 8'h00;
Memory[25649] = 8'h00;
Memory[25648] = 8'h00;
Memory[25655] = 8'h00;
Memory[25654] = 8'h00;
Memory[25653] = 8'h00;
Memory[25652] = 8'h00;
Memory[25659] = 8'h00;
Memory[25658] = 8'h00;
Memory[25657] = 8'h00;
Memory[25656] = 8'h00;
Memory[25663] = 8'h00;
Memory[25662] = 8'h00;
Memory[25661] = 8'h00;
Memory[25660] = 8'h00;
Memory[25667] = 8'h00;
Memory[25666] = 8'h00;
Memory[25665] = 8'h00;
Memory[25664] = 8'h00;
Memory[25671] = 8'h00;
Memory[25670] = 8'h00;
Memory[25669] = 8'h00;
Memory[25668] = 8'h00;
Memory[25675] = 8'h00;
Memory[25674] = 8'h00;
Memory[25673] = 8'h00;
Memory[25672] = 8'h00;
Memory[25679] = 8'h00;
Memory[25678] = 8'h00;
Memory[25677] = 8'h00;
Memory[25676] = 8'h00;
Memory[25683] = 8'h00;
Memory[25682] = 8'h00;
Memory[25681] = 8'h00;
Memory[25680] = 8'h00;
Memory[25687] = 8'h00;
Memory[25686] = 8'h00;
Memory[25685] = 8'h00;
Memory[25684] = 8'h00;
Memory[25691] = 8'h00;
Memory[25690] = 8'h00;
Memory[25689] = 8'h00;
Memory[25688] = 8'h00;
Memory[25695] = 8'h00;
Memory[25694] = 8'h00;
Memory[25693] = 8'h00;
Memory[25692] = 8'h00;
Memory[25699] = 8'h00;
Memory[25698] = 8'h00;
Memory[25697] = 8'h00;
Memory[25696] = 8'h00;
Memory[25703] = 8'h00;
Memory[25702] = 8'h00;
Memory[25701] = 8'h00;
Memory[25700] = 8'h00;
Memory[25707] = 8'h00;
Memory[25706] = 8'h00;
Memory[25705] = 8'h00;
Memory[25704] = 8'h00;
Memory[25711] = 8'h00;
Memory[25710] = 8'h00;
Memory[25709] = 8'h00;
Memory[25708] = 8'h00;
Memory[25715] = 8'h00;
Memory[25714] = 8'h00;
Memory[25713] = 8'h00;
Memory[25712] = 8'h00;
Memory[25719] = 8'h00;
Memory[25718] = 8'h00;
Memory[25717] = 8'h00;
Memory[25716] = 8'h00;
Memory[25723] = 8'h00;
Memory[25722] = 8'h00;
Memory[25721] = 8'h00;
Memory[25720] = 8'h00;
Memory[25727] = 8'h00;
Memory[25726] = 8'h00;
Memory[25725] = 8'h00;
Memory[25724] = 8'h00;
Memory[25731] = 8'h00;
Memory[25730] = 8'h00;
Memory[25729] = 8'h00;
Memory[25728] = 8'h00;
Memory[25735] = 8'h00;
Memory[25734] = 8'h00;
Memory[25733] = 8'h00;
Memory[25732] = 8'h00;
Memory[25739] = 8'h00;
Memory[25738] = 8'h00;
Memory[25737] = 8'h00;
Memory[25736] = 8'h00;
Memory[25743] = 8'h00;
Memory[25742] = 8'h00;
Memory[25741] = 8'h00;
Memory[25740] = 8'h00;
Memory[25747] = 8'h00;
Memory[25746] = 8'h00;
Memory[25745] = 8'h00;
Memory[25744] = 8'h00;
Memory[25751] = 8'h00;
Memory[25750] = 8'h00;
Memory[25749] = 8'h00;
Memory[25748] = 8'h00;
Memory[25755] = 8'h00;
Memory[25754] = 8'h00;
Memory[25753] = 8'h00;
Memory[25752] = 8'h00;
Memory[25759] = 8'h00;
Memory[25758] = 8'h00;
Memory[25757] = 8'h00;
Memory[25756] = 8'h00;
Memory[25763] = 8'h00;
Memory[25762] = 8'h00;
Memory[25761] = 8'h00;
Memory[25760] = 8'h00;
Memory[25767] = 8'h00;
Memory[25766] = 8'h00;
Memory[25765] = 8'h00;
Memory[25764] = 8'h00;
Memory[25771] = 8'h00;
Memory[25770] = 8'h00;
Memory[25769] = 8'h00;
Memory[25768] = 8'h00;
Memory[25775] = 8'h00;
Memory[25774] = 8'h00;
Memory[25773] = 8'h00;
Memory[25772] = 8'h00;
Memory[25779] = 8'h00;
Memory[25778] = 8'h00;
Memory[25777] = 8'h00;
Memory[25776] = 8'h00;
Memory[25783] = 8'h00;
Memory[25782] = 8'h00;
Memory[25781] = 8'h00;
Memory[25780] = 8'h00;
Memory[25787] = 8'h00;
Memory[25786] = 8'h00;
Memory[25785] = 8'h00;
Memory[25784] = 8'h00;
Memory[25791] = 8'h00;
Memory[25790] = 8'h00;
Memory[25789] = 8'h00;
Memory[25788] = 8'h00;
Memory[25795] = 8'h00;
Memory[25794] = 8'h00;
Memory[25793] = 8'h00;
Memory[25792] = 8'h00;
Memory[25799] = 8'h00;
Memory[25798] = 8'h00;
Memory[25797] = 8'h00;
Memory[25796] = 8'h00;
Memory[25803] = 8'h00;
Memory[25802] = 8'h00;
Memory[25801] = 8'h00;
Memory[25800] = 8'h00;
Memory[25807] = 8'h00;
Memory[25806] = 8'h00;
Memory[25805] = 8'h00;
Memory[25804] = 8'h00;
Memory[25811] = 8'h00;
Memory[25810] = 8'h00;
Memory[25809] = 8'h00;
Memory[25808] = 8'h00;
Memory[25815] = 8'h00;
Memory[25814] = 8'h00;
Memory[25813] = 8'h00;
Memory[25812] = 8'h00;
Memory[25819] = 8'h00;
Memory[25818] = 8'h00;
Memory[25817] = 8'h00;
Memory[25816] = 8'h00;
Memory[25823] = 8'h00;
Memory[25822] = 8'h00;
Memory[25821] = 8'h00;
Memory[25820] = 8'h00;
Memory[25827] = 8'h00;
Memory[25826] = 8'h00;
Memory[25825] = 8'h00;
Memory[25824] = 8'h00;
Memory[25831] = 8'h00;
Memory[25830] = 8'h00;
Memory[25829] = 8'h00;
Memory[25828] = 8'h00;
Memory[25835] = 8'h00;
Memory[25834] = 8'h00;
Memory[25833] = 8'h00;
Memory[25832] = 8'h00;
Memory[25839] = 8'h00;
Memory[25838] = 8'h00;
Memory[25837] = 8'h00;
Memory[25836] = 8'h00;
Memory[25843] = 8'h00;
Memory[25842] = 8'h00;
Memory[25841] = 8'h00;
Memory[25840] = 8'h00;
Memory[25847] = 8'h00;
Memory[25846] = 8'h00;
Memory[25845] = 8'h00;
Memory[25844] = 8'h00;
Memory[25851] = 8'h00;
Memory[25850] = 8'h00;
Memory[25849] = 8'h00;
Memory[25848] = 8'h00;
Memory[25855] = 8'h00;
Memory[25854] = 8'h00;
Memory[25853] = 8'h00;
Memory[25852] = 8'h00;
Memory[25859] = 8'h00;
Memory[25858] = 8'h00;
Memory[25857] = 8'h00;
Memory[25856] = 8'h00;
Memory[25863] = 8'h00;
Memory[25862] = 8'h00;
Memory[25861] = 8'h00;
Memory[25860] = 8'h00;
Memory[25867] = 8'h00;
Memory[25866] = 8'h00;
Memory[25865] = 8'h00;
Memory[25864] = 8'h00;
Memory[25871] = 8'h00;
Memory[25870] = 8'h00;
Memory[25869] = 8'h00;
Memory[25868] = 8'h00;
Memory[25875] = 8'h00;
Memory[25874] = 8'h00;
Memory[25873] = 8'h00;
Memory[25872] = 8'h00;
Memory[25879] = 8'h00;
Memory[25878] = 8'h00;
Memory[25877] = 8'h00;
Memory[25876] = 8'h00;
Memory[25883] = 8'h00;
Memory[25882] = 8'h00;
Memory[25881] = 8'h00;
Memory[25880] = 8'h00;
Memory[25887] = 8'h00;
Memory[25886] = 8'h00;
Memory[25885] = 8'h00;
Memory[25884] = 8'h00;
Memory[25891] = 8'h00;
Memory[25890] = 8'h00;
Memory[25889] = 8'h00;
Memory[25888] = 8'h00;
Memory[25895] = 8'h00;
Memory[25894] = 8'h00;
Memory[25893] = 8'h00;
Memory[25892] = 8'h00;
Memory[25899] = 8'h00;
Memory[25898] = 8'h00;
Memory[25897] = 8'h00;
Memory[25896] = 8'h00;
Memory[25903] = 8'h00;
Memory[25902] = 8'h00;
Memory[25901] = 8'h00;
Memory[25900] = 8'h00;
Memory[25907] = 8'h00;
Memory[25906] = 8'h00;
Memory[25905] = 8'h00;
Memory[25904] = 8'h00;
Memory[25911] = 8'h00;
Memory[25910] = 8'h00;
Memory[25909] = 8'h00;
Memory[25908] = 8'h00;
Memory[25915] = 8'h00;
Memory[25914] = 8'h00;
Memory[25913] = 8'h00;
Memory[25912] = 8'h00;
Memory[25919] = 8'h00;
Memory[25918] = 8'h00;
Memory[25917] = 8'h00;
Memory[25916] = 8'h00;
Memory[25923] = 8'h00;
Memory[25922] = 8'h00;
Memory[25921] = 8'h00;
Memory[25920] = 8'h00;
Memory[25927] = 8'h00;
Memory[25926] = 8'h00;
Memory[25925] = 8'h00;
Memory[25924] = 8'h00;
Memory[25931] = 8'h00;
Memory[25930] = 8'h00;
Memory[25929] = 8'h00;
Memory[25928] = 8'h00;
Memory[25935] = 8'h00;
Memory[25934] = 8'h00;
Memory[25933] = 8'h00;
Memory[25932] = 8'h00;
Memory[25939] = 8'h00;
Memory[25938] = 8'h00;
Memory[25937] = 8'h00;
Memory[25936] = 8'h00;
Memory[25943] = 8'h00;
Memory[25942] = 8'h00;
Memory[25941] = 8'h00;
Memory[25940] = 8'h00;
Memory[25947] = 8'h00;
Memory[25946] = 8'h00;
Memory[25945] = 8'h00;
Memory[25944] = 8'h00;
Memory[25951] = 8'h00;
Memory[25950] = 8'h00;
Memory[25949] = 8'h00;
Memory[25948] = 8'h00;
Memory[25955] = 8'h00;
Memory[25954] = 8'h00;
Memory[25953] = 8'h00;
Memory[25952] = 8'h00;
Memory[25959] = 8'h00;
Memory[25958] = 8'h00;
Memory[25957] = 8'h00;
Memory[25956] = 8'h00;
Memory[25963] = 8'h00;
Memory[25962] = 8'h00;
Memory[25961] = 8'h00;
Memory[25960] = 8'h00;
Memory[25967] = 8'h00;
Memory[25966] = 8'h00;
Memory[25965] = 8'h00;
Memory[25964] = 8'h00;
Memory[25971] = 8'h00;
Memory[25970] = 8'h00;
Memory[25969] = 8'h00;
Memory[25968] = 8'h00;
Memory[25975] = 8'h00;
Memory[25974] = 8'h00;
Memory[25973] = 8'h00;
Memory[25972] = 8'h00;
Memory[25979] = 8'h00;
Memory[25978] = 8'h00;
Memory[25977] = 8'h00;
Memory[25976] = 8'h00;
Memory[25983] = 8'h00;
Memory[25982] = 8'h00;
Memory[25981] = 8'h00;
Memory[25980] = 8'h00;
Memory[25987] = 8'h00;
Memory[25986] = 8'h00;
Memory[25985] = 8'h00;
Memory[25984] = 8'h00;
Memory[25991] = 8'h00;
Memory[25990] = 8'h00;
Memory[25989] = 8'h00;
Memory[25988] = 8'h00;
Memory[25995] = 8'h00;
Memory[25994] = 8'h00;
Memory[25993] = 8'h00;
Memory[25992] = 8'h00;
Memory[25999] = 8'h00;
Memory[25998] = 8'h00;
Memory[25997] = 8'h00;
Memory[25996] = 8'h00;
Memory[26003] = 8'h00;
Memory[26002] = 8'h00;
Memory[26001] = 8'h00;
Memory[26000] = 8'h00;
Memory[26007] = 8'h00;
Memory[26006] = 8'h00;
Memory[26005] = 8'h00;
Memory[26004] = 8'h00;
Memory[26011] = 8'h00;
Memory[26010] = 8'h00;
Memory[26009] = 8'h00;
Memory[26008] = 8'h00;
Memory[26015] = 8'h00;
Memory[26014] = 8'h00;
Memory[26013] = 8'h00;
Memory[26012] = 8'h00;
Memory[26019] = 8'h00;
Memory[26018] = 8'h00;
Memory[26017] = 8'h00;
Memory[26016] = 8'h00;
Memory[26023] = 8'h00;
Memory[26022] = 8'h00;
Memory[26021] = 8'h00;
Memory[26020] = 8'h00;
Memory[26027] = 8'h00;
Memory[26026] = 8'h00;
Memory[26025] = 8'h00;
Memory[26024] = 8'h00;
Memory[26031] = 8'h00;
Memory[26030] = 8'h00;
Memory[26029] = 8'h00;
Memory[26028] = 8'h00;
Memory[26035] = 8'h00;
Memory[26034] = 8'h00;
Memory[26033] = 8'h00;
Memory[26032] = 8'h00;
Memory[26039] = 8'h00;
Memory[26038] = 8'h00;
Memory[26037] = 8'h00;
Memory[26036] = 8'h00;
Memory[26043] = 8'h00;
Memory[26042] = 8'h00;
Memory[26041] = 8'h00;
Memory[26040] = 8'h00;
Memory[26047] = 8'h00;
Memory[26046] = 8'h00;
Memory[26045] = 8'h00;
Memory[26044] = 8'h00;
Memory[26051] = 8'h00;
Memory[26050] = 8'h00;
Memory[26049] = 8'h00;
Memory[26048] = 8'h00;
Memory[26055] = 8'h00;
Memory[26054] = 8'h00;
Memory[26053] = 8'h00;
Memory[26052] = 8'h00;
Memory[26059] = 8'h00;
Memory[26058] = 8'h00;
Memory[26057] = 8'h00;
Memory[26056] = 8'h00;
Memory[26063] = 8'h00;
Memory[26062] = 8'h00;
Memory[26061] = 8'h00;
Memory[26060] = 8'h00;
Memory[26067] = 8'h00;
Memory[26066] = 8'h00;
Memory[26065] = 8'h00;
Memory[26064] = 8'h00;
Memory[26071] = 8'h00;
Memory[26070] = 8'h00;
Memory[26069] = 8'h00;
Memory[26068] = 8'h00;
Memory[26075] = 8'h00;
Memory[26074] = 8'h00;
Memory[26073] = 8'h00;
Memory[26072] = 8'h00;
Memory[26079] = 8'h00;
Memory[26078] = 8'h00;
Memory[26077] = 8'h00;
Memory[26076] = 8'h00;
Memory[26083] = 8'h00;
Memory[26082] = 8'h00;
Memory[26081] = 8'h00;
Memory[26080] = 8'h00;
Memory[26087] = 8'h00;
Memory[26086] = 8'h00;
Memory[26085] = 8'h00;
Memory[26084] = 8'h00;
Memory[26091] = 8'h00;
Memory[26090] = 8'h00;
Memory[26089] = 8'h00;
Memory[26088] = 8'h00;
Memory[26095] = 8'h00;
Memory[26094] = 8'h00;
Memory[26093] = 8'h00;
Memory[26092] = 8'h00;
Memory[26099] = 8'h00;
Memory[26098] = 8'h00;
Memory[26097] = 8'h00;
Memory[26096] = 8'h00;
Memory[26103] = 8'h00;
Memory[26102] = 8'h00;
Memory[26101] = 8'h00;
Memory[26100] = 8'h00;
Memory[26107] = 8'h00;
Memory[26106] = 8'h00;
Memory[26105] = 8'h00;
Memory[26104] = 8'h00;
Memory[26111] = 8'h00;
Memory[26110] = 8'h00;
Memory[26109] = 8'h00;
Memory[26108] = 8'h00;
Memory[26115] = 8'h00;
Memory[26114] = 8'h00;
Memory[26113] = 8'h00;
Memory[26112] = 8'h00;
Memory[26119] = 8'h00;
Memory[26118] = 8'h00;
Memory[26117] = 8'h00;
Memory[26116] = 8'h00;
Memory[26123] = 8'h00;
Memory[26122] = 8'h00;
Memory[26121] = 8'h00;
Memory[26120] = 8'h00;
Memory[26127] = 8'h00;
Memory[26126] = 8'h00;
Memory[26125] = 8'h00;
Memory[26124] = 8'h00;
Memory[26131] = 8'h00;
Memory[26130] = 8'h00;
Memory[26129] = 8'h00;
Memory[26128] = 8'h00;
Memory[26135] = 8'h00;
Memory[26134] = 8'h00;
Memory[26133] = 8'h00;
Memory[26132] = 8'h00;
Memory[26139] = 8'h00;
Memory[26138] = 8'h00;
Memory[26137] = 8'h00;
Memory[26136] = 8'h00;
Memory[26143] = 8'h00;
Memory[26142] = 8'h00;
Memory[26141] = 8'h00;
Memory[26140] = 8'h00;
Memory[26147] = 8'h00;
Memory[26146] = 8'h00;
Memory[26145] = 8'h00;
Memory[26144] = 8'h00;
Memory[26151] = 8'h00;
Memory[26150] = 8'h00;
Memory[26149] = 8'h00;
Memory[26148] = 8'h00;
Memory[26155] = 8'h00;
Memory[26154] = 8'h00;
Memory[26153] = 8'h00;
Memory[26152] = 8'h00;
Memory[26159] = 8'h00;
Memory[26158] = 8'h00;
Memory[26157] = 8'h00;
Memory[26156] = 8'h00;
Memory[26163] = 8'h00;
Memory[26162] = 8'h00;
Memory[26161] = 8'h00;
Memory[26160] = 8'h00;
Memory[26167] = 8'h00;
Memory[26166] = 8'h00;
Memory[26165] = 8'h00;
Memory[26164] = 8'h00;
Memory[26171] = 8'h00;
Memory[26170] = 8'h00;
Memory[26169] = 8'h00;
Memory[26168] = 8'h00;
Memory[26175] = 8'h00;
Memory[26174] = 8'h00;
Memory[26173] = 8'h00;
Memory[26172] = 8'h00;
Memory[26179] = 8'h00;
Memory[26178] = 8'h00;
Memory[26177] = 8'h00;
Memory[26176] = 8'h00;
Memory[26183] = 8'h00;
Memory[26182] = 8'h00;
Memory[26181] = 8'h00;
Memory[26180] = 8'h00;
Memory[26187] = 8'h00;
Memory[26186] = 8'h00;
Memory[26185] = 8'h00;
Memory[26184] = 8'h00;
Memory[26191] = 8'h00;
Memory[26190] = 8'h00;
Memory[26189] = 8'h00;
Memory[26188] = 8'h00;
Memory[26195] = 8'h00;
Memory[26194] = 8'h00;
Memory[26193] = 8'h00;
Memory[26192] = 8'h00;
Memory[26199] = 8'h00;
Memory[26198] = 8'h00;
Memory[26197] = 8'h00;
Memory[26196] = 8'h00;
Memory[26203] = 8'h00;
Memory[26202] = 8'h00;
Memory[26201] = 8'h00;
Memory[26200] = 8'h00;
Memory[26207] = 8'h00;
Memory[26206] = 8'h00;
Memory[26205] = 8'h00;
Memory[26204] = 8'h00;
Memory[26211] = 8'h00;
Memory[26210] = 8'h00;
Memory[26209] = 8'h00;
Memory[26208] = 8'h00;
Memory[26215] = 8'h00;
Memory[26214] = 8'h00;
Memory[26213] = 8'h00;
Memory[26212] = 8'h00;
Memory[26219] = 8'h00;
Memory[26218] = 8'h00;
Memory[26217] = 8'h00;
Memory[26216] = 8'h00;
Memory[26223] = 8'h00;
Memory[26222] = 8'h00;
Memory[26221] = 8'h00;
Memory[26220] = 8'h00;
Memory[26227] = 8'h00;
Memory[26226] = 8'h00;
Memory[26225] = 8'h00;
Memory[26224] = 8'h00;
Memory[26231] = 8'h00;
Memory[26230] = 8'h00;
Memory[26229] = 8'h00;
Memory[26228] = 8'h00;
Memory[26235] = 8'h00;
Memory[26234] = 8'h00;
Memory[26233] = 8'h00;
Memory[26232] = 8'h00;
Memory[26239] = 8'h00;
Memory[26238] = 8'h00;
Memory[26237] = 8'h00;
Memory[26236] = 8'h00;
Memory[26243] = 8'h00;
Memory[26242] = 8'h00;
Memory[26241] = 8'h00;
Memory[26240] = 8'h00;
Memory[26247] = 8'h00;
Memory[26246] = 8'h00;
Memory[26245] = 8'h00;
Memory[26244] = 8'h00;
Memory[26251] = 8'h00;
Memory[26250] = 8'h00;
Memory[26249] = 8'h00;
Memory[26248] = 8'h00;
Memory[26255] = 8'h00;
Memory[26254] = 8'h00;
Memory[26253] = 8'h00;
Memory[26252] = 8'h00;
Memory[26259] = 8'h00;
Memory[26258] = 8'h00;
Memory[26257] = 8'h00;
Memory[26256] = 8'h00;

    end
endmodule
