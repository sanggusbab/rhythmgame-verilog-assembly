`timescale  1ns/100ps
module RhythmGameboy_tb();
    reg clk;
    reg[19:0] interrupt;
    wire[7:0] led_A_com;
    wire[7:0] led_A_seg;
    wire[7:0] led_Single;
    wire[11:0] led_RGB;
    wire piezo;
RhythmGameboy RTMGB01(clk, interrupt, led_A_seg, led_A_com, led_Single, led_RGB, piezo);
/*
Reset:      20'b10000000000000000000
Red:        20'b01100000000000000000
Green:      20'b00011000000000000000
Blue:       20'b00000110000000000000
Pause:      20'b00000001000000000000
1key:       20'b00000000100000000000
2key:       20'b00000000010000000000
3key:       20'b00000000001000000000
4key:       20'b00000000000100000000
5key:       20'b00000000000010000000
6key:       20'b00000000000001000000
7key:       20'b00000000000000100000
8key:       20'b00000000000000010000
9key:       20'b00000000000000001000
starkey:    20'b00000000000000000100
0key:       20'b00000000000000000010
hashkey:    20'b00000000000000000001
*/
    always begin
        #5 clk = ~clk;
    end
    initial begin
        interrupt = 20'b0;
        clk = 0;
        #30000 interrupt = 20'b00100000000000000000;
        #30000 interrupt = 20'b01000000000000000000;
        #30000 interrupt = 20'b01100000000000000000;
        #30000 interrupt = 20'b00011000000000000000;
        #30000 interrupt = 20'b00000110000000000000;
        #30000 interrupt = 20'b01111110000000000000;
        #30000 interrupt = 20'b00000000000000000001; // Status 1
        #30000 interrupt = 20'b00000000000000000000;
        #30000 interrupt = 20'b00000000000000000001; // Status 2
        #30000 interrupt = 20'b00000000000000000000;
        #30000 interrupt = 20'b00000000000000010000; // Status 3
        #30000 interrupt = 20'b00000000000000000000;
        #30000 interrupt = 20'b00000000000000010000; // Status 4
        #30000 interrupt = 20'b00000000000000000000;
        #30000 interrupt = 20'b00000000000000010000; // Status 5
        #30000 interrupt = 20'b00000000000000000000;
        #30000 interrupt = 20'b00000000000000000100; // Status 8
        #30000 interrupt = 20'b00000000000000000000;
        #30000 interrupt = 20'b00000000000001000000; // Status 9
        #30000 interrupt = 20'b00000000000000000000;
        #30000 interrupt = 20'b00000000000000000100; // Status 10
        #30000 interrupt = 20'b00000000000000000000;
        #30000 interrupt = 20'b00000000000001000000; // Status 11
        #30000 interrupt = 20'b00000000000000000000;
        #30000 interrupt = 20'b00000000000001000000; // Status 12
        #30000 interrupt = 20'b00000000000000000000;
        #30000 interrupt = 20'b00000000000001000000; // Status 13
        #30000 interrupt = 20'b00000000000000000000;
        #30000 interrupt = 20'b00000000000100000000; // Status 12
        #30000 interrupt = 20'b00000000000000000000;
        #30000 interrupt = 20'b00000000000000000001; // Status 9
        #30000 interrupt = 20'b00000000000000000000;
        #30000 interrupt = 20'b00000000000001000000; // Status 19
        #30000 interrupt = 20'b00000000000000000000;
        #30000 interrupt = 20'b00000000000000000100; // Status 20
        #30000 interrupt = 20'b00000000000000000000;
        #30000 interrupt = 20'b00000000000001000000; // Status 21
        #30000 interrupt = 20'b00000000000000000000;
        #30000 interrupt = 20'b00000000000001000000; // Status 22
        #30000 interrupt = 20'b00000000000000000000;
        #30000 interrupt = 20'b00000000000001000000; // Status 23
        #30000 interrupt = 20'b00000000000000000000;
        #30000 interrupt = 20'b00000000000001000000; // Status 24
        #30000 interrupt = 20'b00000000000000000000;
        #30000 interrupt = 20'b00000000000001000000; // Status 25
        #30000 interrupt = 20'b00000000000000000000;
        #30000 interrupt = 20'b00000000000001000000; // Status 26
        #30000 interrupt = 20'b00000000000000000000;
        #30000 interrupt = 20'b00000000000001000000; // Status 27
        #30000 interrupt = 20'b00000000000000000000;
        #30000 interrupt = 20'b00000000000000000001; // Status 19
        #30000 interrupt = 20'b00000000000000000000;
        #30000 interrupt = 20'b00000000000001000000; // Status 28
        #30000 interrupt = 20'b00000000000000000000;
        #30000 interrupt = 20'b00000000000000000100; // Status 29
        #30000 interrupt = 20'b00000000000000000000;
        #30000 interrupt = 20'b00000000000000000100; // Status 30
        #30000 interrupt = 20'b00000000000000000000;
        #30000 interrupt = 20'b00000000010000000000;
        #30000 interrupt = 20'b00000000000000000000;
        #30000 interrupt = 20'b00000000100000000000;
        #30000 interrupt = 20'b00000000000000000000;
        #30000 interrupt = 20'b00000000000000000010; // 210
        #30000 interrupt = 20'b00000000000000000000;
        #30000 interrupt = 20'b00000000000000000100; // Status 29
        #30000 interrupt = 20'b00000000000000000000;
        #30000 interrupt = 20'b00000000000000010000; // Status 31
        #30000 interrupt = 20'b00000000000000000000;
        #30000 interrupt = 20'b00000000000000000100; // Status 32
        #30000 interrupt = 20'b00000000000000000000;
        #30000 interrupt = 20'b00000000000000000001; // Status 31
        #30000 interrupt = 20'b00000000000000000000;
        #30000 interrupt = 20'b00000000000000000001; // Status 33
        #30000 interrupt = 20'b00000000000000000000;
        #30000 interrupt = 20'b00000000000100000000; // Status 19
        #30000 interrupt = 20'b00000000000000000000;
        #30000 interrupt = 20'b00000000000100000000; // Status 9
        #30000 interrupt = 20'b00000000000000000000;
        #30000 interrupt = 20'b00000000000100000000; // Status 8
        #30000 interrupt = 20'b00000000000000000000;
        #30000 interrupt = 20'b00000000000000000100; // Status 37
        #30000 interrupt = 20'b00000000000000000000;
        #30000 interrupt = 20'b00000000000001000000; // Status 38
        #30000 interrupt = 20'b00000000000000000000;
        #30000 interrupt = 20'b00000000000100000000; // Status 37
        #30000 interrupt = 20'b00000000000000000000;
        #30000 interrupt = 20'b00000000000000000100; // Status 41
        #30000 interrupt = 20'b00000000000000000000;
        #30000 interrupt = 20'b00000000000000010000; // Status 42
        #30000 interrupt = 20'b00000000000000000000;
        #30000 interrupt = 20'b00000000010000000000; // Status 41
        #30000 interrupt = 20'b00000000000000000000;
        #30000 interrupt = 20'b00000000000000000100; // Status 43
        #30000 interrupt = 20'b00000000000000000000;
        #1000000000;
        #1000000000;
        #1000000000;
        #1000000000;
        #1000000000 interrupt = 20'b00000001000000000000; // Status 46
        #30000 interrupt = 20'b00000001000000010000; // Status 49
        #30000 interrupt = 20'b00000001000000000000;
        #30000 interrupt = 20'b00000001010000000000; // Status 46
        #30000 interrupt = 20'b00000001000000000000;
        #30000 interrupt = 20'b00000001010000000000; // Status 48
        #30000 interrupt = 20'b00000001000000000000;
        #30000 interrupt = 20'b00000001010000000000; // Status 47
        #30000 interrupt = 20'b00000001000000000000;
        #30000 interrupt = 20'b00000001000000000100; // Status 50
        #30000 interrupt = 20'b00000001000000000000;
        #30000 interrupt = 20'b00000001000000000100; // Status 43
        #30000 interrupt = 20'b00000001000000000000;
        #30000 interrupt = 20'b00000000000000000000;
    end
endmodule
